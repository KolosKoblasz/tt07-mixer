magic
tech sky130A
magscale 1 2
timestamp 1716477521
<< pwell >>
rect -201 -717 201 717
<< psubdiff >>
rect -165 647 -69 681
rect 69 647 165 681
rect -165 585 -131 647
rect 131 585 165 647
rect -165 -647 -131 -585
rect 131 -647 165 -585
rect -165 -681 -69 -647
rect 69 -681 165 -647
<< psubdiffcont >>
rect -69 647 69 681
rect -165 -585 -131 585
rect 131 -585 165 585
rect -69 -681 69 -647
<< xpolycontact >>
rect -35 119 35 551
rect -35 -551 35 -119
<< xpolyres >>
rect -35 -119 35 119
<< locali >>
rect -165 647 -69 681
rect 69 647 165 681
rect -165 585 -131 647
rect 131 585 165 647
rect -165 -647 -131 -585
rect 131 -647 165 -585
rect -165 -681 -69 -647
rect 69 -681 165 -647
<< viali >>
rect -19 136 19 533
rect -19 -533 19 -136
<< metal1 >>
rect -25 533 25 545
rect -25 136 -19 533
rect 19 136 25 533
rect -25 124 25 136
rect -25 -136 25 -124
rect -25 -533 -19 -136
rect 19 -533 25 -136
rect -25 -545 25 -533
<< properties >>
string FIXED_BBOX -148 -664 148 664
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.35 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 8.789k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
