magic
tech sky130A
magscale 1 2
timestamp 1716477521
<< locali >>
rect -100 250 100 307
rect -100 -307 100 -250
<< rlocali >>
rect -100 -250 100 250
<< properties >>
string gencell sky130_fd_pr__res_generic_l1
string library sky130
string parameters w 1 l 2.5 m 1 nx 1 wmin 0.17 lmin 0.17 rho 12.8 val 32.0 dummy 0 dw 0.0 term 0.0 snake 0 roverlap 0
<< end >>
