magic
tech sky130A
magscale 1 2
timestamp 1716477521
<< locali >>
rect -40 100 40 157
rect -40 -157 40 -100
<< rlocali >>
rect -40 -100 40 100
<< properties >>
string gencell sky130_fd_pr__res_generic_l1
string library sky130
string parameters w 0.4 l 1 m 1 nx 1 wmin 0.17 lmin 0.17 rho 12.8 val 32.0 dummy 0 dw 0.0 term 0.0 snake 0 roverlap 0
<< end >>
