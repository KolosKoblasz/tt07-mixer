magic
tech sky130A
magscale 1 2
timestamp 1717082701
<< metal1 >>
rect 28190 19800 28200 20200
rect 28400 19800 30000 20200
rect 28190 19000 28200 19400
rect 28400 19000 29200 19400
rect 28800 18400 29200 19000
rect 29600 18400 30000 19800
rect 24790 17600 24800 18000
rect 25000 17600 27000 18000
rect 26990 16400 27000 16800
rect 27200 16400 27400 16800
rect 31190 16400 31200 16800
rect 31400 16400 31410 16800
rect 25990 15400 26000 15600
rect 26400 15400 27800 15600
rect 26000 15200 27800 15400
rect 30800 15400 32000 15600
rect 32400 15400 32410 15600
rect 30800 15200 32400 15400
rect 24790 14200 24800 14600
rect 25000 14200 29400 14600
<< via1 >>
rect 28200 19800 28400 20200
rect 28200 19000 28400 19400
rect 24800 17600 25000 18000
rect 27000 16400 27200 16800
rect 31200 16400 31400 16800
rect 26000 15400 26400 15600
rect 32000 15400 32400 15600
rect 24800 14200 25000 14600
<< metal2 >>
rect 25800 43100 25900 43110
rect 12100 43000 25800 43100
rect 12100 41400 12200 43000
rect 25800 42990 25900 43000
rect 26600 42900 26700 42910
rect 14000 42800 26600 42900
rect 14000 41400 14100 42800
rect 26600 42790 26700 42800
rect 27300 42700 27400 42710
rect 15900 42600 27300 42700
rect 15900 41400 16100 42600
rect 27300 42590 27400 42600
rect 28000 42500 28100 42510
rect 17900 42400 28000 42500
rect 17900 41400 18000 42400
rect 28000 42390 28100 42400
rect 28800 42300 28900 42310
rect 19800 42200 28800 42300
rect 19800 41400 19900 42200
rect 28800 42190 28900 42200
rect 29500 42100 29600 42110
rect 21700 42000 29500 42100
rect 21700 41400 21900 42000
rect 29500 41990 29600 42000
rect 30200 41900 30300 41910
rect 23700 41800 30200 41900
rect 23700 41400 23800 41800
rect 30200 41790 30300 41800
rect 30949 41667 31056 41671
rect 25624 41662 31061 41667
rect 25624 41555 30949 41662
rect 31056 41555 31061 41662
rect 25624 41550 31061 41555
rect 25624 41396 25680 41550
rect 30949 41546 31056 41550
rect 27600 37400 27800 37410
rect 27800 37000 30000 37400
rect 27600 36990 27800 37000
rect 27400 29400 27600 29410
rect 27600 29000 29200 29400
rect 27400 28990 27600 29000
rect 28800 21200 29200 29000
rect 26000 20800 29200 21200
rect 29600 21200 30000 37000
rect 29600 20800 32400 21200
rect 24000 18400 24200 18410
rect 24200 18000 25000 18400
rect 24200 17600 24800 18000
rect 24000 17590 24200 17600
rect 24800 17590 25000 17600
rect 26000 15600 26400 20800
rect 27600 20200 27800 20210
rect 28200 20200 28400 20210
rect 27800 19800 28200 20200
rect 27600 19790 27800 19800
rect 28200 19790 28400 19800
rect 27600 19400 27800 19410
rect 28200 19400 28400 19410
rect 27800 19000 28200 19400
rect 27600 18990 27800 19000
rect 28200 18990 28400 19000
rect 27000 16800 27200 16810
rect 26800 16400 27000 16800
rect 26800 16000 27200 16400
rect 26800 15790 27200 15800
rect 31200 16800 31400 16810
rect 31400 16400 31600 16800
rect 31200 16000 31600 16400
rect 31200 15790 31600 15800
rect 26000 15390 26400 15400
rect 32000 15600 32400 20800
rect 32000 15390 32400 15400
rect 24000 14800 24200 14810
rect 24200 14600 25000 14800
rect 24200 14200 24800 14600
rect 24200 14000 25000 14200
rect 24000 13990 24200 14000
<< via2 >>
rect 25800 43000 25900 43100
rect 26600 42800 26700 42900
rect 27300 42600 27400 42700
rect 28000 42400 28100 42500
rect 28800 42200 28900 42300
rect 29500 42000 29600 42100
rect 30200 41800 30300 41900
rect 30949 41555 31056 41662
rect 27600 37000 27800 37400
rect 27400 29000 27600 29400
rect 24000 17600 24200 18400
rect 27600 19800 27800 20200
rect 27600 19000 27800 19400
rect 26800 15800 27200 16000
rect 31200 15800 31600 16000
rect 24000 14000 24200 14800
<< metal3 >>
rect 25790 44900 25800 45000
rect 25900 44900 25910 45000
rect 26590 44900 26600 45000
rect 26700 44900 26710 45000
rect 27290 44900 27300 45000
rect 27400 44900 27410 45000
rect 27990 44900 28000 45000
rect 28100 44900 28110 45000
rect 28790 44900 28800 45000
rect 28900 44900 28910 45000
rect 29490 44900 29500 45000
rect 29600 44900 29610 45000
rect 30190 44900 30200 45000
rect 30300 44900 30310 45000
rect 30950 44932 31062 44938
rect 30950 44908 30960 44932
rect 25800 43105 25900 44900
rect 25790 43100 25910 43105
rect 25790 43000 25800 43100
rect 25900 43000 25910 43100
rect 25790 42995 25910 43000
rect 26600 42905 26700 44900
rect 26590 42900 26710 42905
rect 26590 42800 26600 42900
rect 26700 42800 26710 42900
rect 26590 42795 26710 42800
rect 27300 42705 27400 44900
rect 27290 42700 27410 42705
rect 27290 42600 27300 42700
rect 27400 42600 27410 42700
rect 27290 42595 27410 42600
rect 28000 42505 28100 44900
rect 27990 42500 28110 42505
rect 27990 42400 28000 42500
rect 28100 42400 28110 42500
rect 27990 42395 28110 42400
rect 28800 42305 28900 44900
rect 28790 42300 28910 42305
rect 28790 42200 28800 42300
rect 28900 42200 28910 42300
rect 28790 42195 28910 42200
rect 29500 42105 29600 44900
rect 29490 42100 29610 42105
rect 29490 42000 29500 42100
rect 29600 42000 29610 42100
rect 29490 41995 29610 42000
rect 30200 41905 30300 44900
rect 30944 44866 30960 44908
rect 31050 44866 31062 44932
rect 30944 44832 31062 44866
rect 30190 41900 30310 41905
rect 30190 41800 30200 41900
rect 30300 41800 30310 41900
rect 30190 41795 30310 41800
rect 30944 41662 31061 44832
rect 30944 41555 30949 41662
rect 31056 41555 31061 41662
rect 30944 41550 31061 41555
rect 27590 37400 27810 37405
rect 26800 37000 27600 37400
rect 27800 37000 27810 37400
rect 27590 36995 27810 37000
rect 27390 29400 27610 29405
rect 26600 29000 27400 29400
rect 27600 29000 27610 29400
rect 27390 28995 27610 29000
rect 13126 24946 13426 24952
rect 20552 24946 20852 24952
rect 201 24328 499 24333
rect 13126 24328 13426 24646
rect 16810 24934 17110 24946
rect 16810 24328 17110 24634
rect 20552 24328 20852 24646
rect 24236 24946 24536 24952
rect 24236 24328 24536 24646
rect 200 24327 24536 24328
rect 200 24029 201 24327
rect 499 24029 24536 24327
rect 200 24028 24536 24029
rect 201 24023 499 24028
rect 27590 20200 27810 20205
rect 26990 19800 27000 20200
rect 27200 19800 27600 20200
rect 27800 19800 27810 20200
rect 27590 19795 27810 19800
rect 27590 19400 27810 19405
rect 26990 19000 27000 19400
rect 27200 19000 27600 19400
rect 27800 19000 27810 19400
rect 27590 18995 27810 19000
rect 1990 17400 2000 18600
rect 2200 18405 24200 18600
rect 2200 18400 24210 18405
rect 2200 17600 24000 18400
rect 24200 17600 24210 18400
rect 2200 17595 24210 17600
rect 2200 17400 24200 17595
rect 26790 16000 27210 16005
rect 26790 15800 26800 16000
rect 27200 15800 27210 16000
rect 26790 15795 27210 15800
rect 31190 16000 31610 16005
rect 31190 15800 31200 16000
rect 31600 15800 31610 16000
rect 31190 15795 31610 15800
rect 26800 15600 27200 15795
rect 31200 15600 31600 15795
rect 26790 15400 26800 15600
rect 27200 15400 27210 15600
rect 31190 15400 31200 15600
rect 31600 15400 31610 15600
rect 11990 13800 12000 15000
rect 12200 14805 24200 15000
rect 12200 14800 24210 14805
rect 12200 14000 24000 14800
rect 24200 14000 24210 14800
rect 12200 13995 24210 14000
rect 12200 13800 24200 13995
<< via3 >>
rect 25800 44900 25900 45000
rect 26600 44900 26700 45000
rect 27300 44900 27400 45000
rect 28000 44900 28100 45000
rect 28800 44900 28900 45000
rect 29500 44900 29600 45000
rect 30200 44900 30300 45000
rect 30960 44866 31050 44932
rect 13126 24646 13426 24946
rect 16810 24634 17110 24934
rect 20552 24646 20852 24946
rect 24236 24646 24536 24946
rect 201 24029 499 24327
rect 27000 19800 27200 20200
rect 27000 19000 27200 19400
rect 2000 17400 2200 18600
rect 26800 15400 27200 15600
rect 31200 15400 31600 15600
rect 12000 13800 12200 15000
<< metal4 >>
rect 798 45000 858 45152
rect 1534 45000 1594 45152
rect 2270 45000 2330 45152
rect 3006 45000 3066 45152
rect 3742 45000 3802 45152
rect 4478 45000 4538 45152
rect 5214 45000 5274 45152
rect 5950 45000 6010 45152
rect 6686 45000 6746 45152
rect 7422 45000 7482 45152
rect 8158 45000 8218 45152
rect 8894 45000 8954 45152
rect 9630 45000 9690 45152
rect 10366 45000 10426 45152
rect 11102 45000 11162 45152
rect 11838 45000 11898 45152
rect 12574 45000 12634 45152
rect 13310 45000 13370 45152
rect 14046 45000 14106 45152
rect 14782 45000 14842 45152
rect 15518 45000 15578 45152
rect 16254 45000 16314 45152
rect 16990 45000 17050 45152
rect 17726 45000 17786 45152
rect 600 44800 17800 45000
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44950 24410 45152
rect 25086 44952 25146 45152
rect 25822 45001 25882 45152
rect 26558 45001 26618 45152
rect 27294 45001 27354 45152
rect 28030 45001 28090 45152
rect 28766 45001 28826 45152
rect 29502 45001 29562 45152
rect 30238 45002 30298 45152
rect 30196 45001 30300 45002
rect 25799 45000 25901 45001
rect 26558 45000 26701 45001
rect 27294 45000 27401 45001
rect 25799 44900 25800 45000
rect 25900 44900 25901 45000
rect 26500 44900 26600 45000
rect 26700 44900 26701 45000
rect 27200 44900 27300 45000
rect 27400 44900 27401 45000
rect 25799 44899 25901 44900
rect 26599 44899 26701 44900
rect 27299 44899 27401 44900
rect 27999 45000 28101 45001
rect 28766 45000 28901 45001
rect 27999 44900 28000 45000
rect 28100 44900 28101 45000
rect 28700 44900 28800 45000
rect 28900 44900 28901 45000
rect 27999 44899 28101 44900
rect 28799 44899 28901 44900
rect 29499 45000 29601 45001
rect 29499 44900 29500 45000
rect 29600 44900 29601 45000
rect 29499 44899 29601 44900
rect 30196 45000 30301 45001
rect 30196 44900 30200 45000
rect 30300 44900 30301 45000
rect 30974 44939 31034 45152
rect 31710 44952 31770 45152
rect 30196 44899 30301 44900
rect 30953 44932 31063 44939
rect 30196 44896 30300 44899
rect 30953 44866 30960 44932
rect 31050 44866 31063 44932
rect 30953 44857 31063 44866
rect 9800 44552 10200 44800
rect 9790 44460 10200 44552
rect 200 24327 500 44152
rect 9790 43994 10194 44460
rect 200 24029 201 24327
rect 499 24029 500 24327
rect 200 18600 500 24029
rect 1999 18600 2201 18601
rect 200 17400 2000 18600
rect 2200 17400 2201 18600
rect 200 1000 500 17400
rect 1999 17399 2201 17400
rect 9800 15086 10100 43994
rect 13126 24947 13426 26206
rect 13125 24946 13427 24947
rect 13125 24646 13126 24946
rect 13426 24646 13427 24946
rect 13125 24645 13427 24646
rect 14990 23750 15290 26204
rect 16810 24935 17110 26162
rect 16809 24934 17111 24935
rect 16809 24634 16810 24934
rect 17110 24634 17111 24934
rect 16809 24633 17111 24634
rect 18690 23750 18990 26126
rect 20552 24947 20852 26226
rect 20551 24946 20853 24947
rect 20551 24646 20552 24946
rect 20852 24646 20853 24946
rect 20551 24645 20853 24646
rect 22386 23750 22686 26148
rect 24236 24947 24536 26130
rect 26082 25702 26382 26194
rect 26064 25528 26382 25702
rect 24235 24946 24537 24947
rect 24235 24646 24236 24946
rect 24536 24646 24537 24946
rect 24235 24645 24537 24646
rect 26064 23750 26364 25528
rect 10292 23450 26364 23750
rect 22386 23448 22686 23450
rect 26999 20200 27201 20201
rect 19800 19800 27000 20200
rect 27200 19800 27201 20200
rect 9800 15000 10466 15086
rect 11999 15000 12201 15001
rect 9800 13800 12000 15000
rect 12200 13800 12201 15000
rect 9800 13644 10466 13800
rect 11999 13799 12201 13800
rect 9800 1000 10100 13644
rect 19800 3200 20200 19800
rect 26999 19799 27201 19800
rect 26999 19400 27201 19401
rect 18000 2800 20200 3200
rect 20600 19000 27000 19400
rect 27200 19000 27201 19400
rect 20600 3200 21000 19000
rect 26999 18999 27201 19000
rect 26799 15600 27201 15601
rect 26799 15400 26800 15600
rect 27200 15400 27201 15600
rect 26799 15399 27201 15400
rect 31199 15600 31601 15601
rect 31199 15400 31200 15600
rect 31600 15400 31601 15600
rect 31199 15399 31601 15400
rect 26800 13400 27200 15399
rect 31200 13400 31600 15399
rect 26800 13000 29000 13400
rect 28600 3200 29000 13000
rect 20600 2800 22800 3200
rect 18000 430 18400 2800
rect 22400 430 22800 2800
rect 26800 2800 29000 3200
rect 29400 13000 31600 13400
rect 29400 3200 29800 13000
rect 29400 2800 31600 3200
rect 26800 434 27200 2800
rect 31200 434 31600 2800
rect 26864 432 27200 434
rect 31280 432 31600 434
rect 18032 276 18214 430
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 276
rect 22450 0 22630 430
rect 26866 0 27046 432
rect 31282 430 31600 432
rect 31282 0 31462 430
use gilbert_mixer  gilbert_mixer_0
timestamp 1716553577
transform 1 0 26624 0 1 16514
box 200 -2000 4600 2000
use mixer_control  mixer_control_0
timestamp 1717082701
transform 1 0 10886 0 1 25468
box 514 496 16000 16000
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
