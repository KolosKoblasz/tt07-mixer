* NGSPICE file created from gilbert_mixer_parax.ext - technology: sky130A

.subckt gilbert_mixer_parax VSS VDD OUT_N OUT_P LO_N LO_P IN_N IN_P
X0 OUT_N.t0 VDD.t0 VSS.t0 sky130_fd_pr__res_xhigh_po_0p35 l=1.35
X1 NET_M6_DRAIN IN_P.t0 OUT_N.t1 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=0.38
X2 NET_M5_DRAIN IN_P.t1 OUT_P.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=0.38
X3 NET_M5_DRAIN IN_N.t0 OUT_N.t3 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=0.38
X4 OUT_N.t4 IN_P.t2 NET_M6_DRAIN VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=0.38
X5 OUT_P.t4 IN_N.t1 NET_M6_DRAIN VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=0.38
X6 OUT_N.t2 IN_N.t2 NET_M5_DRAIN VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=0.38
X7 NET_M6_DRAIN IN_N.t3 OUT_P.t3 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=0.38
X8 VDD.t1 OUT_P.t2 VSS.t7 sky130_fd_pr__res_xhigh_po_0p35 l=1.35
X9 NET_R3 LO_P.t0 NET_M5_DRAIN VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=0.38
R0 NET_R3 VSS sky130_fd_pr__res_generic_l1 w=0.4 l=1
X10 NET_M5_DRAIN LO_P.t1 NET_R3 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=0.38
X11 NET_R3 LO_N.t0 NET_M6_DRAIN VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=0.38
X12 NET_M6_DRAIN LO_N.t1 NET_R3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=0.38
X13 OUT_P.t0 IN_P.t3 NET_M5_DRAIN VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=0.38
R1 OUT_N.n1 OUT_N.t4 51.1305
R2 OUT_N.n0 OUT_N.t3 51.1305
R3 OUT_N.n1 OUT_N.t1 50.9487
R4 OUT_N.n0 OUT_N.t2 50.9487
R5 OUT_N.n3 OUT_N.t0 42.5533
R6 OUT_N OUT_N.n3 2.973
R7 OUT_N.n3 OUT_N.n2 1.5357
R8 OUT_N.n2 OUT_N.n0 0.176971
R9 OUT_N.n2 OUT_N.n1 0.176971
R10 VDD.n0 VDD.t0 43.8786
R11 VDD.n0 VDD.t1 42.5516
R12 VDD.n1 VDD.n0 0.437132
R13 VDD.n1 VDD 0.0702115
R14 VDD VDD.n1 0.0688962
R15 VSS.n83 VSS.n12 4606.32
R16 VSS.n71 VSS.n12 4606.32
R17 VSS.n83 VSS.n13 4606.32
R18 VSS.n71 VSS.n13 4606.32
R19 VSS.n56 VSS.n18 4606.32
R20 VSS.n56 VSS.n19 4606.32
R21 VSS.n57 VSS.n18 4606.32
R22 VSS.n57 VSS.n19 4606.32
R23 VSS.n74 VSS.n62 3291.06
R24 VSS.n74 VSS.n63 3291.06
R25 VSS.n70 VSS.n62 3291.06
R26 VSS.n70 VSS.n63 3291.06
R27 VSS.n86 VSS.n6 3291.06
R28 VSS.n90 VSS.n6 3291.06
R29 VSS.n86 VSS.n7 3291.06
R30 VSS.n90 VSS.n7 3291.06
R31 VSS.n45 VSS.n24 3291.06
R32 VSS.n45 VSS.n25 3291.06
R33 VSS.n24 VSS.n23 3291.06
R34 VSS.n25 VSS.n23 3291.06
R35 VSS.n93 VSS.n4 3291.06
R36 VSS.n67 VSS.n4 3291.06
R37 VSS.n93 VSS.n5 3291.06
R38 VSS.n67 VSS.n5 3291.06
R39 VSS.n53 VSS.n21 3291.06
R40 VSS.n53 VSS.n48 3291.06
R41 VSS.n21 VSS.n20 3291.06
R42 VSS.n48 VSS.n20 3291.06
R43 VSS.n33 VSS.n30 3291.06
R44 VSS.n38 VSS.n30 3291.06
R45 VSS.n33 VSS.n31 3291.06
R46 VSS.n38 VSS.n31 3291.06
R47 VSS.n85 VSS.n10 554.4
R48 VSS.n72 VSS.n71 512.5
R49 VSS.n34 VSS.n18 327.7
R50 VSS.n82 VSS.n14 299.295
R51 VSS.n15 VSS.n14 299.295
R52 VSS.n82 VSS.n81 299.295
R53 VSS.n55 VSS.n16 299.295
R54 VSS.n55 VSS.n17 299.295
R55 VSS.n58 VSS.n17 299.295
R56 VSS.n19 VSS.n17 292.5
R57 VSS.n19 VSS.n10 292.5
R58 VSS.n18 VSS.n16 292.5
R59 VSS.n71 VSS.n15 292.5
R60 VSS.n83 VSS.n82 292.5
R61 VSS.n84 VSS.n83 292.5
R62 VSS.n69 VSS.n61 213.835
R63 VSS.n69 VSS.n60 213.835
R64 VSS.n88 VSS.n87 213.835
R65 VSS.n89 VSS.n88 213.835
R66 VSS.n44 VSS.n26 213.835
R67 VSS.n44 VSS.n43 213.835
R68 VSS.n66 VSS.n2 213.835
R69 VSS.n66 VSS.n3 213.835
R70 VSS.n94 VSS.n3 213.835
R71 VSS.n52 VSS.n51 213.835
R72 VSS.n51 VSS.n50 213.835
R73 VSS.n50 VSS.n49 213.835
R74 VSS.n39 VSS.n29 213.835
R75 VSS.n32 VSS.n29 213.835
R76 VSS.t10 VSS.n34 199.101
R77 VSS.t3 VSS.n10 199.101
R78 VSS.t4 VSS.n72 199.101
R79 VSS.n59 VSS.n16 196.769
R80 VSS.n27 VSS.n26 195.886
R81 VSS.n32 VSS.n28 195.886
R82 VSS.n75 VSS.n61 195.644
R83 VSS.n89 VSS.n8 195.644
R84 VSS.n43 VSS.n42 195.388
R85 VSS.n40 VSS.n39 195.388
R86 VSS.n76 VSS.n60 193.656
R87 VSS.n87 VSS.n9 193.656
R88 VSS.n85 VSS.n84 184.8
R89 VSS.n80 VSS.n15 163.341
R90 VSS.n52 VSS.n1 143.963
R91 VSS.n95 VSS.n2 140.549
R92 VSS.n50 VSS.n20 117.001
R93 VSS.n54 VSS.n20 117.001
R94 VSS.n53 VSS.n52 117.001
R95 VSS.n54 VSS.n53 117.001
R96 VSS.n5 VSS.n3 117.001
R97 VSS.n64 VSS.n5 117.001
R98 VSS.n4 VSS.n2 117.001
R99 VSS.n64 VSS.n4 117.001
R100 VSS.n27 VSS.n23 117.001
R101 VSS.n46 VSS.n23 117.001
R102 VSS.n45 VSS.n44 117.001
R103 VSS.n46 VSS.n45 117.001
R104 VSS.n88 VSS.n7 117.001
R105 VSS.n11 VSS.n7 117.001
R106 VSS.n8 VSS.n6 117.001
R107 VSS.n11 VSS.n6 117.001
R108 VSS.n70 VSS.n69 117.001
R109 VSS.n73 VSS.n70 117.001
R110 VSS.n75 VSS.n74 117.001
R111 VSS.n74 VSS.n73 117.001
R112 VSS.n30 VSS.n29 117.001
R113 VSS.n35 VSS.n30 117.001
R114 VSS.n31 VSS.n28 117.001
R115 VSS.n35 VSS.n31 117.001
R116 VSS.n37 VSS.n36 105.6
R117 VSS.n47 VSS.n22 105.6
R118 VSS.n92 VSS.n91 105.6
R119 VSS.n36 VSS.t8 93.5005
R120 VSS.n37 VSS.t2 93.5005
R121 VSS.n22 VSS.t1 93.5005
R122 VSS.n47 VSS.t12 93.5005
R123 VSS.n92 VSS.t11 93.5005
R124 VSS.n91 VSS.t5 93.5005
R125 VSS.n65 VSS.t6 93.5005
R126 VSS.t13 VSS.n68 93.5005
R127 VSS.n35 VSS.t10 73.7005
R128 VSS.t8 VSS.n35 73.7005
R129 VSS.n54 VSS.t1 73.7005
R130 VSS.t12 VSS.n46 73.7005
R131 VSS.n46 VSS.t3 73.7005
R132 VSS.t9 VSS.n11 73.7005
R133 VSS.n11 VSS.t11 73.7005
R134 VSS.n64 VSS.t5 73.7005
R135 VSS.t6 VSS.n64 73.7005
R136 VSS.n73 VSS.t13 73.7005
R137 VSS.n73 VSS.t4 73.7005
R138 VSS.n49 VSS.n48 73.1255
R139 VSS.n48 VSS.n47 73.1255
R140 VSS.n51 VSS.n21 73.1255
R141 VSS.n36 VSS.n21 73.1255
R142 VSS.n67 VSS.n66 73.1255
R143 VSS.n68 VSS.n67 73.1255
R144 VSS.n94 VSS.n93 73.1255
R145 VSS.n93 VSS.n92 73.1255
R146 VSS.n43 VSS.n25 73.1255
R147 VSS.n25 VSS.n10 73.1255
R148 VSS.n26 VSS.n24 73.1255
R149 VSS.n24 VSS.n22 73.1255
R150 VSS.n90 VSS.n89 73.1255
R151 VSS.n91 VSS.n90 73.1255
R152 VSS.n87 VSS.n86 73.1255
R153 VSS.n86 VSS.n85 73.1255
R154 VSS.n63 VSS.n61 73.1255
R155 VSS.n72 VSS.n63 73.1255
R156 VSS.n62 VSS.n60 73.1255
R157 VSS.n65 VSS.n62 73.1255
R158 VSS.n39 VSS.n38 73.1255
R159 VSS.n38 VSS.n37 73.1255
R160 VSS.n33 VSS.n32 73.1255
R161 VSS.n34 VSS.n33 73.1255
R162 VSS.n68 VSS.t7 70.4005
R163 VSS.n81 VSS.n80 68.8476
R164 VSS.t0 VSS.t2 56.1005
R165 VSS.n49 VSS.n1 50.5981
R166 VSS.n59 VSS.n58 50.3221
R167 VSS.n95 VSS.n94 47.1848
R168 VSS.t7 VSS.n65 35.2005
R169 VSS.n58 VSS.n57 34.4123
R170 VSS.n57 VSS.t0 34.4123
R171 VSS.n56 VSS.n55 34.4123
R172 VSS.t0 VSS.n56 34.4123
R173 VSS.n81 VSS.n13 34.4123
R174 VSS.t7 VSS.n13 34.4123
R175 VSS.n14 VSS.n12 34.4123
R176 VSS.t7 VSS.n12 34.4123
R177 VSS.t0 VSS.n54 17.6005
R178 VSS.n84 VSS.t9 14.3005
R179 VSS.n78 VSS.n77 8.39189
R180 VSS.n41 VSS.n0 8.13618
R181 VSS.n96 VSS.n1 5.05362
R182 VSS.n96 VSS.n95 5.0505
R183 VSS.n80 VSS.n79 4.62672
R184 VSS.n79 VSS.n59 4.5104
R185 VSS.n77 VSS.n76 3.5755
R186 VSS.n41 VSS.n40 2.9505
R187 VSS.n97 VSS.n96 2.8305
R188 VSS.n77 VSS.n9 2.3255
R189 VSS.n42 VSS.n41 2.3255
R190 VSS VSS.n97 2.22873
R191 VSS.n76 VSS.n75 1.0245
R192 VSS.n9 VSS.n8 1.0245
R193 VSS.n42 VSS.n27 0.2565
R194 VSS.n40 VSS.n28 0.2565
R195 VSS.n78 VSS.n0 0.17619
R196 VSS.n97 VSS.n0 0.138143
R197 VSS.n79 VSS.n78 0.0900238
R198 IN_P.n4 IN_P.t3 310.603
R199 IN_P.t2 IN_P.n1 310.579
R200 IN_P.n2 IN_P.t2 310.579
R201 IN_P.t3 IN_P.n0 310.579
R202 IN_P.n2 IN_P.t0 310.339
R203 IN_P.t0 IN_P.n1 310.339
R204 IN_P.t1 IN_P.n0 310.339
R205 IN_P.n4 IN_P.t1 310.339
R206 IN_P.n5 IN_P.n3 3.53502
R207 IN_P.n3 IN_P.n1 1.32014
R208 IN_P.n5 IN_P.n4 0.588
R209 IN_P.n6 IN_P.n0 0.588
R210 IN_P.n3 IN_P.n2 0.570143
R211 IN_P.n6 IN_P.n5 0.393357
R212 IN_P IN_P.n6 0.191125
R213 OUT_P.n0 OUT_P.t3 50.9487
R214 OUT_P.n1 OUT_P.t1 50.9372
R215 OUT_P.n0 OUT_P.t4 50.9357
R216 OUT_P.n1 OUT_P.t0 50.9106
R217 OUT_P.n2 OUT_P.t2 43.2255
R218 OUT_P OUT_P.n3 2.14737
R219 OUT_P.n3 OUT_P.n0 1.3408
R220 OUT_P.n2 OUT_P.n1 0.502732
R221 OUT_P.n3 OUT_P.n2 0.340344
R222 IN_N.n4 IN_N.t3 310.579
R223 IN_N.n1 IN_N.t0 310.579
R224 IN_N.t0 IN_N.n0 310.579
R225 IN_N.n5 IN_N.t3 310.579
R226 IN_N.n1 IN_N.t2 310.339
R227 IN_N.t2 IN_N.n0 310.339
R228 IN_N.t1 IN_N.n4 310.339
R229 IN_N.n5 IN_N.t1 310.339
R230 IN_N.n3 IN_N.n2 12.8392
R231 IN_N.n2 IN_N.n0 1.3136
R232 IN_N IN_N.n5 0.638
R233 IN_N.n4 IN_N.n3 0.504071
R234 IN_N.n2 IN_N.n1 0.464389
R235 IN_N IN_N.n3 0.354667
R236 LO_P.n1 LO_P.t1 310.579
R237 LO_P.t1 LO_P.n0 310.579
R238 LO_P.t0 LO_P.n0 310.339
R239 LO_P.n1 LO_P.t0 310.339
R240 LO_P.n2 LO_P.n1 1.01955
R241 LO_P.n2 LO_P.n0 0.561214
R242 LO_P LO_P.n2 0.2005
R243 LO_N.t0 LO_N.n0 310.579
R244 LO_N.n1 LO_N.t0 310.579
R245 LO_N.t1 LO_N.n0 310.339
R246 LO_N.n1 LO_N.t1 310.339
R247 LO_N LO_N.n0 1.03383
R248 LO_N LO_N.n1 0.649029
C0 LO_N LO_P 0.002325f
C1 OUT_P LO_N 4.08e-19
C2 NET_M5_DRAIN LO_P 0.38819f
C3 OUT_P NET_M5_DRAIN 0.706311f
C4 OUT_N LO_N 5.83e-21
C5 OUT_N NET_M5_DRAIN 0.659731f
C6 LO_N NET_M6_DRAIN 0.386256f
C7 OUT_P VDD 0.480519f
C8 OUT_P LO_P 4.06e-19
C9 NET_R3 li_2560_n1733# 0.021591f
C10 NET_M6_DRAIN NET_M5_DRAIN 0.011342f
C11 NET_R3 IN_P 0.00259f
C12 OUT_N VDD 0.468992f
C13 OUT_P OUT_N 1.20018f
C14 IN_N NET_R3 0.008931f
C15 NET_M6_DRAIN VDD 2.21e-19
C16 NET_M6_DRAIN LO_P 3.45e-21
C17 OUT_P NET_M6_DRAIN 0.69523f
C18 OUT_N NET_M6_DRAIN 0.671935f
C19 IN_N IN_P 0.566608f
C20 LO_N NET_R3 0.166236f
C21 NET_M5_DRAIN NET_R3 0.707667f
C22 NET_R3 LO_P 0.170642f
C23 NET_M5_DRAIN IN_P 0.340914f
C24 OUT_N NET_R3 0.020856f
C25 LO_N IN_N 0.094715f
C26 NET_M5_DRAIN IN_N 0.20055f
C27 NET_M6_DRAIN NET_R3 0.69861f
C28 VDD IN_P 0.035515f
C29 LO_P IN_P 0.074279f
C30 OUT_P IN_P 0.412796f
C31 OUT_N IN_P 0.654526f
C32 IN_N VDD 0.015363f
C33 OUT_P IN_N 0.484173f
C34 NET_M6_DRAIN IN_P 0.17147f
C35 OUT_N IN_N 0.571687f
C36 NET_M6_DRAIN IN_N 0.353623f
C37 LO_N NET_M5_DRAIN 3.45e-21
C38 LO_N VSS 1.16427f
C39 LO_P VSS 1.18326f
C40 IN_N VSS 3.80717f
C41 IN_P VSS 3.12094f
C42 OUT_N VSS 3.31039f
C43 OUT_P VSS 5.1178f
C44 VDD VSS 3.72634f
C45 li_2560_n1733# VSS 0.139933f $ **FLOATING
C46 NET_R3 VSS 1.47547f
C47 NET_M6_DRAIN VSS 1.38852f
C48 NET_M5_DRAIN VSS 1.14576f
.ends

