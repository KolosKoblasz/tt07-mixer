magic
tech sky130A
magscale 1 2
timestamp 1716482002
<< viali >>
rect 1090 810 1400 890
rect 3560 820 3880 880
rect 1150 320 1460 360
rect 1950 320 2260 360
rect 2950 -380 3250 -330
rect 3750 -380 4050 -330
rect 1930 -1130 1990 -970
rect 3220 -1130 3270 -970
rect 2580 -1530 2620 -1490
rect 2580 -1780 2620 -1740
<< metal1 >>
rect 2200 1970 2400 2000
rect 2200 1820 2230 1970
rect 2360 1820 2400 1970
rect 2200 1800 2400 1820
rect 3000 1800 3200 2000
rect 200 1404 934 1408
rect 200 1400 3800 1404
rect 200 1200 4080 1400
rect 320 1196 4080 1200
rect 910 1190 1440 1196
rect 960 940 1400 1190
rect 3010 1050 3020 1060
rect 1070 890 1420 900
rect 1070 810 1090 890
rect 1400 810 1420 890
rect 1070 770 1420 810
rect 1640 680 2070 1040
rect 1640 590 1660 680
rect 2060 590 2070 680
rect 1640 580 2070 590
rect 2950 930 3020 1050
rect 3180 1050 3190 1060
rect 3180 930 3400 1050
rect 3600 940 4080 1196
rect 2950 490 3400 930
rect 3540 880 3900 900
rect 3540 820 3560 880
rect 3880 820 3900 880
rect 3540 800 3900 820
rect 2950 410 2960 490
rect 3380 410 3400 490
rect 2340 380 2440 400
rect 2950 390 3400 410
rect 1120 360 2360 380
rect 1120 320 1150 360
rect 1460 320 1950 360
rect 2260 320 2360 360
rect 2420 320 2440 380
rect 1120 300 2440 320
rect 870 200 1410 270
rect 1970 200 2510 270
rect 600 0 940 200
rect 1130 0 1140 170
rect 1200 0 1210 170
rect 1390 0 1400 170
rect 1480 0 1490 170
rect 1920 10 1930 160
rect 2000 10 2010 160
rect 2190 10 2200 160
rect 2260 10 2270 160
rect 870 -220 940 0
rect 1260 -170 1270 -60
rect 1330 -170 1340 -60
rect 2060 -170 2070 -60
rect 2130 -170 2140 -60
rect 2440 -170 2510 200
rect 2420 -210 2510 -170
rect 2420 -220 2440 -210
rect 870 -230 1240 -220
rect 870 -290 1410 -230
rect 1960 -280 2440 -220
rect 2500 -280 2510 -210
rect 1960 -290 2510 -280
rect 2680 200 3220 270
rect 3780 200 4320 270
rect 2680 -220 2750 200
rect 2930 10 2940 160
rect 3000 10 3010 160
rect 3190 10 3200 160
rect 3270 10 3280 160
rect 3730 10 3740 160
rect 3800 10 3810 160
rect 3990 10 4000 160
rect 4070 10 4080 160
rect 4250 0 4600 200
rect 3060 -180 3070 -50
rect 3140 -180 3150 -50
rect 3860 -180 3870 -50
rect 3930 -180 3940 -50
rect 4250 -220 4340 0
rect 2680 -290 3220 -220
rect 3770 -290 4340 -220
rect 870 -435 940 -290
rect 2680 -435 2750 -290
rect 870 -510 2750 -435
rect 2930 -330 4100 -320
rect 2930 -380 2950 -330
rect 3250 -380 3750 -330
rect 4050 -380 4100 -330
rect 2930 -400 4100 -380
rect 2930 -470 2960 -400
rect 3070 -470 4100 -400
rect 2930 -480 4100 -470
rect 4250 -540 4340 -290
rect 2430 -550 4340 -540
rect 2500 -610 4340 -550
rect 2430 -620 4340 -610
rect 1290 -1000 1820 -930
rect 1920 -970 3290 -950
rect 1000 -1200 1350 -1000
rect 1530 -1180 1540 -1040
rect 1600 -1180 1610 -1040
rect 1800 -1180 1810 -1040
rect 1870 -1180 1880 -1040
rect 1920 -1130 1930 -970
rect 1990 -990 3220 -970
rect 1990 -1110 2530 -990
rect 2670 -1110 3220 -990
rect 1990 -1130 3220 -1110
rect 3270 -1130 3290 -970
rect 3390 -1000 3920 -930
rect 1920 -1150 3290 -1130
rect 3330 -1180 3340 -1050
rect 3400 -1180 3410 -1050
rect 3600 -1180 3610 -1050
rect 3670 -1180 3680 -1050
rect 1290 -1420 1350 -1200
rect 3860 -1200 4200 -1000
rect 2530 -1240 2670 -1230
rect 1660 -1380 1670 -1240
rect 1730 -1380 1740 -1240
rect 2530 -1370 2540 -1240
rect 2660 -1370 2670 -1240
rect 3460 -1370 3470 -1240
rect 3530 -1370 3540 -1240
rect 1290 -1490 1820 -1420
rect 2530 -1490 2670 -1370
rect 3860 -1420 3920 -1200
rect 3390 -1490 3920 -1420
rect 2530 -1530 2580 -1490
rect 2620 -1530 2670 -1490
rect 2530 -1550 2670 -1530
rect 2540 -1740 2670 -1660
rect 2540 -1780 2580 -1740
rect 2620 -1780 2670 -1740
rect 2540 -1800 2670 -1780
rect 2500 -1830 2700 -1800
rect 2500 -1980 2530 -1830
rect 2670 -1980 2700 -1830
rect 2500 -2000 2700 -1980
<< via1 >>
rect 2230 1820 2360 1970
rect 1090 810 1400 890
rect 1660 590 2060 680
rect 3020 930 3180 1060
rect 3560 820 3880 880
rect 2960 410 3380 490
rect 2360 320 2420 380
rect 1140 0 1200 170
rect 1400 0 1480 170
rect 1930 10 2000 160
rect 2200 10 2260 160
rect 1270 -170 1330 -60
rect 2070 -170 2130 -60
rect 2440 -280 2500 -210
rect 2940 10 3000 160
rect 3200 10 3270 160
rect 3740 10 3800 160
rect 4000 10 4070 160
rect 3070 -180 3140 -50
rect 3870 -180 3930 -50
rect 2960 -470 3070 -400
rect 2430 -610 2500 -550
rect 1540 -1180 1600 -1040
rect 1810 -1180 1870 -1040
rect 2530 -1110 2670 -990
rect 3340 -1180 3400 -1050
rect 3610 -1180 3670 -1050
rect 1670 -1380 1730 -1240
rect 2540 -1370 2660 -1240
rect 3470 -1370 3530 -1240
rect 2530 -1980 2670 -1830
<< metal2 >>
rect 2220 1970 2370 1980
rect 2220 1820 2230 1970
rect 2360 1820 2370 1970
rect 1070 890 1420 900
rect 1070 810 1090 890
rect 1400 810 1420 890
rect 1070 770 1420 810
rect 2220 740 2370 1820
rect 3010 1060 3180 1990
rect 3010 930 3020 1060
rect 3010 920 3180 930
rect 3540 880 3900 900
rect 3540 820 3560 880
rect 3880 820 3900 880
rect 3540 800 3900 820
rect 1130 680 4080 740
rect 1130 590 1660 680
rect 2060 590 4080 680
rect 1130 580 4080 590
rect 1130 170 1480 580
rect 2470 490 3400 510
rect 2470 410 2960 490
rect 3380 410 3400 490
rect 2340 380 2440 400
rect 2340 320 2360 380
rect 2420 320 2440 380
rect 2340 300 2440 320
rect 2470 390 3400 410
rect 2470 170 2730 390
rect 1130 0 1140 170
rect 1200 0 1400 170
rect 1930 160 3270 170
rect 2000 10 2200 160
rect 2260 10 2940 160
rect 3000 10 3200 160
rect 1930 0 3270 10
rect 3740 160 4080 580
rect 3800 10 4000 160
rect 4070 10 4080 160
rect 3740 0 4080 10
rect 1140 -10 1200 0
rect 1400 -10 1480 0
rect 3070 -50 3140 -40
rect 3870 -50 3930 -40
rect 1260 -60 2140 -50
rect 1260 -170 1270 -60
rect 1330 -170 2070 -60
rect 2130 -170 2140 -60
rect 1260 -180 2140 -170
rect 3140 -180 3870 -50
rect 3930 -180 3950 -50
rect 1630 -1040 1800 -180
rect 3070 -190 3140 -180
rect 2430 -210 2500 -200
rect 2430 -280 2440 -210
rect 2430 -550 2500 -280
rect 2920 -400 3100 -390
rect 2920 -470 2960 -400
rect 3070 -470 3100 -400
rect 2920 -480 3100 -470
rect 2430 -620 2500 -610
rect 2510 -990 2690 -970
rect 1520 -1180 1540 -1040
rect 1600 -1180 1810 -1040
rect 1870 -1180 1890 -1040
rect 2510 -1110 2530 -990
rect 2670 -1110 2690 -990
rect 3410 -1040 3580 -180
rect 3870 -190 3930 -180
rect 2510 -1130 2690 -1110
rect 3320 -1050 3690 -1040
rect 1520 -1190 1890 -1180
rect 3320 -1180 3340 -1050
rect 3400 -1180 3610 -1050
rect 3670 -1180 3690 -1050
rect 3320 -1190 3690 -1180
rect 1660 -1240 3540 -1230
rect 1660 -1380 1670 -1240
rect 1730 -1370 2540 -1240
rect 2660 -1370 3470 -1240
rect 3530 -1370 3540 -1240
rect 1730 -1380 3540 -1370
rect 1670 -1390 1730 -1380
rect 2500 -1830 2700 -1800
rect 2500 -1980 2530 -1830
rect 2670 -1980 2700 -1830
rect 2500 -2000 2700 -1980
<< via2 >>
rect 1090 810 1400 890
rect 3560 820 3880 880
rect 2360 320 2420 380
rect 2960 -470 3070 -400
rect 2530 -1110 2670 -990
rect 2530 -1980 2670 -1830
<< metal3 >>
rect 1070 890 1420 900
rect 1070 810 1090 890
rect 1400 810 1420 890
rect 1070 800 1420 810
rect 3540 880 3900 900
rect 3540 820 3560 880
rect 3880 820 3900 880
rect 3540 800 3900 820
rect 1070 700 3900 800
rect 2500 400 2710 700
rect 2340 380 2710 400
rect 2340 320 2360 380
rect 2420 320 2710 380
rect 2340 300 2710 320
rect 2500 -390 2710 300
rect 2500 -400 3100 -390
rect 2500 -470 2960 -400
rect 3070 -470 3100 -400
rect 2500 -480 3100 -470
rect 2500 -990 2710 -480
rect 2500 -1110 2530 -990
rect 2670 -1110 2710 -990
rect 2500 -1830 2710 -1110
rect 2500 -1980 2530 -1830
rect 2670 -1980 2710 -1830
rect 2500 -2000 2710 -1980
use sky130_fd_pr__res_generic_l1_TPAW2P  sky130_fd_pr__res_generic_l1_TPAW2P_0
timestamp 1716477521
transform 1 0 2600 0 1 -1633
box -40 -157 40 157
use sky130_fd_pr__res_xhigh_po_0p35_EFWLNN  sky130_fd_pr__res_xhigh_po_0p35_EFWLNN_0
timestamp 1716477521
transform 0 1 3517 -1 0 1001
box -201 -717 201 717
use sky130_fd_pr__res_xhigh_po_0p35_EFWLNN  sky130_fd_pr__res_xhigh_po_0p35_EFWLNN_1
timestamp 1716477521
transform 0 1 1517 -1 0 1001
box -201 -717 201 717
use sky130_fd_pr__nfet_01v8_WX3E3J  XM1 ~/projects/tt07-mixer/mag
timestamp 1716455288
transform 1 0 2101 0 1 -10
box -301 -390 301 390
use sky130_fd_pr__nfet_01v8_WX3E3J  XM2
timestamp 1716455288
transform 1 0 1701 0 1 -1210
box -301 -390 301 390
use sky130_fd_pr__nfet_01v8_WX3E3J  XM3
timestamp 1716455288
transform 1 0 3101 0 1 -10
box -301 -390 301 390
use sky130_fd_pr__nfet_01v8_WX3E3J  XM4
timestamp 1716455288
transform 1 0 3501 0 1 -1210
box -301 -390 301 390
use sky130_fd_pr__nfet_01v8_WX3E3J  XM5
timestamp 1716455288
transform 1 0 3901 0 1 -10
box -301 -390 301 390
use sky130_fd_pr__nfet_01v8_WX3E3J  XM6
timestamp 1716455288
transform 1 0 1301 0 1 -10
box -301 -390 301 390
<< labels >>
flabel metal1 4000 -1200 4200 -1000 0 FreeSans 256 0 0 0 LO_N
port 4 nsew
flabel metal1 1000 -1200 1200 -1000 0 FreeSans 256 0 0 0 LO_P
port 5 nsew
flabel metal1 600 0 800 200 0 FreeSans 256 0 0 0 IN_P
port 7 nsew
flabel metal1 2200 1800 2400 2000 0 FreeSans 256 0 0 0 OUT_P
port 3 nsew
flabel metal1 4400 0 4600 200 0 FreeSans 256 0 0 0 IN_N
port 6 nsew
flabel metal2 1630 -1190 1800 -50 0 FreeSans 480 0 0 0 NET_M5_DRAIN
flabel metal2 3410 -1190 3580 -50 0 FreeSans 480 0 0 0 NET_M6_DRAIN
flabel metal1 3000 1800 3200 2000 0 FreeSans 256 0 0 0 OUT_N
port 2 nsew
flabel metal1 204 1204 404 1404 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel via1 2540 -1370 2660 -1240 0 FreeSans 480 0 0 0 NET_R3
flabel metal1 2500 -2000 2700 -1800 0 FreeSans 256 0 0 0 VSS
port 0 nsew
<< end >>
