magic
tech sky130A
magscale 1 2
timestamp 1716477521
<< pwell >>
rect -685 -761 685 761
<< psubdiff >>
rect -649 691 -553 725
rect 553 691 649 725
rect -649 629 -615 691
rect 615 629 649 691
rect -649 -691 -615 -629
rect 615 -691 649 -629
rect -649 -725 -553 -691
rect 553 -725 649 -691
<< psubdiffcont >>
rect -553 691 553 725
rect -649 -629 -615 629
rect 615 -629 649 629
rect -553 -725 553 -691
<< poly >>
rect -519 579 -453 595
rect -519 545 -503 579
rect -469 545 -453 579
rect -519 165 -453 545
rect -519 -545 -453 -165
rect -519 -579 -503 -545
rect -469 -579 -453 -545
rect -519 -595 -453 -579
rect -411 579 -345 595
rect -411 545 -395 579
rect -361 545 -345 579
rect -411 165 -345 545
rect -411 -545 -345 -165
rect -411 -579 -395 -545
rect -361 -579 -345 -545
rect -411 -595 -345 -579
rect -303 579 -237 595
rect -303 545 -287 579
rect -253 545 -237 579
rect -303 165 -237 545
rect -303 -545 -237 -165
rect -303 -579 -287 -545
rect -253 -579 -237 -545
rect -303 -595 -237 -579
rect -195 579 -129 595
rect -195 545 -179 579
rect -145 545 -129 579
rect -195 165 -129 545
rect -195 -545 -129 -165
rect -195 -579 -179 -545
rect -145 -579 -129 -545
rect -195 -595 -129 -579
rect -87 579 -21 595
rect -87 545 -71 579
rect -37 545 -21 579
rect -87 165 -21 545
rect -87 -545 -21 -165
rect -87 -579 -71 -545
rect -37 -579 -21 -545
rect -87 -595 -21 -579
rect 21 579 87 595
rect 21 545 37 579
rect 71 545 87 579
rect 21 165 87 545
rect 21 -545 87 -165
rect 21 -579 37 -545
rect 71 -579 87 -545
rect 21 -595 87 -579
rect 129 579 195 595
rect 129 545 145 579
rect 179 545 195 579
rect 129 165 195 545
rect 129 -545 195 -165
rect 129 -579 145 -545
rect 179 -579 195 -545
rect 129 -595 195 -579
rect 237 579 303 595
rect 237 545 253 579
rect 287 545 303 579
rect 237 165 303 545
rect 237 -545 303 -165
rect 237 -579 253 -545
rect 287 -579 303 -545
rect 237 -595 303 -579
rect 345 579 411 595
rect 345 545 361 579
rect 395 545 411 579
rect 345 165 411 545
rect 345 -545 411 -165
rect 345 -579 361 -545
rect 395 -579 411 -545
rect 345 -595 411 -579
rect 453 579 519 595
rect 453 545 469 579
rect 503 545 519 579
rect 453 165 519 545
rect 453 -545 519 -165
rect 453 -579 469 -545
rect 503 -579 519 -545
rect 453 -595 519 -579
<< polycont >>
rect -503 545 -469 579
rect -503 -579 -469 -545
rect -395 545 -361 579
rect -395 -579 -361 -545
rect -287 545 -253 579
rect -287 -579 -253 -545
rect -179 545 -145 579
rect -179 -579 -145 -545
rect -71 545 -37 579
rect -71 -579 -37 -545
rect 37 545 71 579
rect 37 -579 71 -545
rect 145 545 179 579
rect 145 -579 179 -545
rect 253 545 287 579
rect 253 -579 287 -545
rect 361 545 395 579
rect 361 -579 395 -545
rect 469 545 503 579
rect 469 -579 503 -545
<< npolyres >>
rect -519 -165 -453 165
rect -411 -165 -345 165
rect -303 -165 -237 165
rect -195 -165 -129 165
rect -87 -165 -21 165
rect 21 -165 87 165
rect 129 -165 195 165
rect 237 -165 303 165
rect 345 -165 411 165
rect 453 -165 519 165
<< locali >>
rect -649 691 -553 725
rect 553 691 649 725
rect -649 629 -615 691
rect 615 629 649 691
rect -519 545 -503 579
rect -469 545 -453 579
rect -411 545 -395 579
rect -361 545 -345 579
rect -303 545 -287 579
rect -253 545 -237 579
rect -195 545 -179 579
rect -145 545 -129 579
rect -87 545 -71 579
rect -37 545 -21 579
rect 21 545 37 579
rect 71 545 87 579
rect 129 545 145 579
rect 179 545 195 579
rect 237 545 253 579
rect 287 545 303 579
rect 345 545 361 579
rect 395 545 411 579
rect 453 545 469 579
rect 503 545 519 579
rect -519 -579 -503 -545
rect -469 -579 -453 -545
rect -411 -579 -395 -545
rect -361 -579 -345 -545
rect -303 -579 -287 -545
rect -253 -579 -237 -545
rect -195 -579 -179 -545
rect -145 -579 -129 -545
rect -87 -579 -71 -545
rect -37 -579 -21 -545
rect 21 -579 37 -545
rect 71 -579 87 -545
rect 129 -579 145 -545
rect 179 -579 195 -545
rect 237 -579 253 -545
rect 287 -579 303 -545
rect 345 -579 361 -545
rect 395 -579 411 -545
rect 453 -579 469 -545
rect 503 -579 519 -545
rect -649 -691 -615 -629
rect 615 -691 649 -629
rect -649 -725 -553 -691
rect 553 -725 649 -691
<< viali >>
rect -503 545 -469 579
rect -395 545 -361 579
rect -287 545 -253 579
rect -179 545 -145 579
rect -71 545 -37 579
rect 37 545 71 579
rect 145 545 179 579
rect 253 545 287 579
rect 361 545 395 579
rect 469 545 503 579
rect -503 182 -469 545
rect -395 182 -361 545
rect -287 182 -253 545
rect -179 182 -145 545
rect -71 182 -37 545
rect 37 182 71 545
rect 145 182 179 545
rect 253 182 287 545
rect 361 182 395 545
rect 469 182 503 545
rect -503 -545 -469 -182
rect -395 -545 -361 -182
rect -287 -545 -253 -182
rect -179 -545 -145 -182
rect -71 -545 -37 -182
rect 37 -545 71 -182
rect 145 -545 179 -182
rect 253 -545 287 -182
rect 361 -545 395 -182
rect 469 -545 503 -182
rect -503 -579 -469 -545
rect -395 -579 -361 -545
rect -287 -579 -253 -545
rect -179 -579 -145 -545
rect -71 -579 -37 -545
rect 37 -579 71 -545
rect 145 -579 179 -545
rect 253 -579 287 -545
rect 361 -579 395 -545
rect 469 -579 503 -545
<< metal1 >>
rect -509 579 -463 591
rect -509 182 -503 579
rect -469 182 -463 579
rect -509 170 -463 182
rect -401 579 -355 591
rect -401 182 -395 579
rect -361 182 -355 579
rect -401 170 -355 182
rect -293 579 -247 591
rect -293 182 -287 579
rect -253 182 -247 579
rect -293 170 -247 182
rect -185 579 -139 591
rect -185 182 -179 579
rect -145 182 -139 579
rect -185 170 -139 182
rect -77 579 -31 591
rect -77 182 -71 579
rect -37 182 -31 579
rect -77 170 -31 182
rect 31 579 77 591
rect 31 182 37 579
rect 71 182 77 579
rect 31 170 77 182
rect 139 579 185 591
rect 139 182 145 579
rect 179 182 185 579
rect 139 170 185 182
rect 247 579 293 591
rect 247 182 253 579
rect 287 182 293 579
rect 247 170 293 182
rect 355 579 401 591
rect 355 182 361 579
rect 395 182 401 579
rect 355 170 401 182
rect 463 579 509 591
rect 463 182 469 579
rect 503 182 509 579
rect 463 170 509 182
rect -509 -182 -463 -170
rect -509 -579 -503 -182
rect -469 -579 -463 -182
rect -509 -591 -463 -579
rect -401 -182 -355 -170
rect -401 -579 -395 -182
rect -361 -579 -355 -182
rect -401 -591 -355 -579
rect -293 -182 -247 -170
rect -293 -579 -287 -182
rect -253 -579 -247 -182
rect -293 -591 -247 -579
rect -185 -182 -139 -170
rect -185 -579 -179 -182
rect -145 -579 -139 -182
rect -185 -591 -139 -579
rect -77 -182 -31 -170
rect -77 -579 -71 -182
rect -37 -579 -31 -182
rect -77 -591 -31 -579
rect 31 -182 77 -170
rect 31 -579 37 -182
rect 71 -579 77 -182
rect 31 -591 77 -579
rect 139 -182 185 -170
rect 139 -579 145 -182
rect 179 -579 185 -182
rect 139 -591 185 -579
rect 247 -182 293 -170
rect 247 -579 253 -182
rect 287 -579 293 -182
rect 247 -591 293 -579
rect 355 -182 401 -170
rect 355 -579 361 -182
rect 395 -579 401 -182
rect 355 -591 401 -579
rect 463 -182 509 -170
rect 463 -579 469 -182
rect 503 -579 509 -182
rect 463 -591 509 -579
<< properties >>
string FIXED_BBOX -632 -708 632 708
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.330 l 1.650 m 1 nx 10 wmin 0.330 lmin 1.650 rho 48.2 val 241.0 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
