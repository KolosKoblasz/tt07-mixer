magic
tech sky130A
magscale 1 2
timestamp 1716901194
<< viali >>
rect 9413 15113 9447 15147
rect 4353 15045 4387 15079
rect 7389 15045 7423 15079
rect 3525 14977 3559 15011
rect 4169 14977 4203 15011
rect 10977 14977 11011 15011
rect 1317 14909 1351 14943
rect 3341 14909 3375 14943
rect 4445 14909 4479 14943
rect 5181 14909 5215 14943
rect 6377 14909 6411 14943
rect 6469 14909 6503 14943
rect 7021 14909 7055 14943
rect 7205 14909 7239 14943
rect 8585 14909 8619 14943
rect 8861 14909 8895 14943
rect 9229 14909 9263 14943
rect 9689 14909 9723 14943
rect 11253 14909 11287 14943
rect 12909 14909 12943 14943
rect 1501 14773 1535 14807
rect 4445 14773 4479 14807
rect 5365 14773 5399 14807
rect 6285 14773 6319 14807
rect 8769 14773 8803 14807
rect 9045 14773 9079 14807
rect 10333 14773 10367 14807
rect 11897 14773 11931 14807
rect 13093 14773 13127 14807
rect 4813 14569 4847 14603
rect 9505 14569 9539 14603
rect 9597 14569 9631 14603
rect 5273 14501 5307 14535
rect 5825 14501 5859 14535
rect 14105 14501 14139 14535
rect 3709 14433 3743 14467
rect 4169 14433 4203 14467
rect 4353 14433 4387 14467
rect 4445 14433 4479 14467
rect 4629 14433 4663 14467
rect 5089 14433 5123 14467
rect 5365 14433 5399 14467
rect 5457 14433 5491 14467
rect 6101 14433 6135 14467
rect 7409 14433 7443 14467
rect 7665 14433 7699 14467
rect 7757 14433 7791 14467
rect 8024 14433 8058 14467
rect 10241 14433 10275 14467
rect 11437 14433 11471 14467
rect 14013 14433 14047 14467
rect 3617 14365 3651 14399
rect 4077 14365 4111 14399
rect 5825 14365 5859 14399
rect 9413 14365 9447 14399
rect 11713 14365 11747 14399
rect 13185 14365 13219 14399
rect 13829 14365 13863 14399
rect 4537 14297 4571 14331
rect 5641 14297 5675 14331
rect 6285 14297 6319 14331
rect 9137 14297 9171 14331
rect 9965 14297 9999 14331
rect 6009 14229 6043 14263
rect 10149 14229 10183 14263
rect 13277 14229 13311 14263
rect 4721 14025 4755 14059
rect 5641 14025 5675 14059
rect 7665 14025 7699 14059
rect 8401 14025 8435 14059
rect 11897 14025 11931 14059
rect 12725 14025 12759 14059
rect 4353 13957 4387 13991
rect 6837 13957 6871 13991
rect 6193 13889 6227 13923
rect 6285 13889 6319 13923
rect 7021 13889 7055 13923
rect 7849 13889 7883 13923
rect 9137 13889 9171 13923
rect 12357 13889 12391 13923
rect 12449 13889 12483 13923
rect 4261 13821 4295 13855
rect 4537 13821 4571 13855
rect 5822 13821 5856 13855
rect 6561 13821 6595 13855
rect 6653 13821 6687 13855
rect 7757 13821 7791 13855
rect 7941 13821 7975 13855
rect 8585 13821 8619 13855
rect 8861 13821 8895 13855
rect 9045 13821 9079 13855
rect 9321 13821 9355 13855
rect 9413 13821 9447 13855
rect 9597 13821 9631 13855
rect 9689 13821 9723 13855
rect 11805 13821 11839 13855
rect 12725 13821 12759 13855
rect 12909 13821 12943 13855
rect 13001 13821 13035 13855
rect 13737 13821 13771 13855
rect 6837 13753 6871 13787
rect 5825 13685 5859 13719
rect 10333 13685 10367 13719
rect 12265 13685 12299 13719
rect 13185 13685 13219 13719
rect 13553 13685 13587 13719
rect 4721 13481 4755 13515
rect 10333 13481 10367 13515
rect 7573 13413 7607 13447
rect 10977 13413 11011 13447
rect 5089 13345 5123 13379
rect 7665 13345 7699 13379
rect 10149 13345 10183 13379
rect 10425 13345 10459 13379
rect 10609 13345 10643 13379
rect 5181 13277 5215 13311
rect 5273 13277 5307 13311
rect 9965 13277 9999 13311
rect 10517 13277 10551 13311
rect 6285 13141 6319 13175
rect 7849 13141 7883 13175
rect 12265 13141 12299 13175
rect 4813 12937 4847 12971
rect 5457 12937 5491 12971
rect 5641 12937 5675 12971
rect 6745 12937 6779 12971
rect 10977 12937 11011 12971
rect 5089 12801 5123 12835
rect 5181 12733 5215 12767
rect 5917 12733 5951 12767
rect 6653 12733 6687 12767
rect 8125 12733 8159 12767
rect 9781 12733 9815 12767
rect 12357 12733 12391 12767
rect 6285 12665 6319 12699
rect 6469 12665 6503 12699
rect 7858 12665 7892 12699
rect 9514 12665 9548 12699
rect 12112 12665 12146 12699
rect 8401 12597 8435 12631
rect 5365 12393 5399 12427
rect 7021 12393 7055 12427
rect 7205 12393 7239 12427
rect 9137 12393 9171 12427
rect 9321 12393 9355 12427
rect 4905 12257 4939 12291
rect 8493 12257 8527 12291
rect 9229 12257 9263 12291
rect 9413 12257 9447 12291
rect 14565 12257 14599 12291
rect 6653 12189 6687 12223
rect 5181 12053 5215 12087
rect 7021 12053 7055 12087
rect 14749 12053 14783 12087
rect 11345 4709 11379 4743
rect 11253 4437 11287 4471
<< metal1 >>
rect 552 15258 15364 15280
rect 552 15206 2249 15258
rect 2301 15206 2313 15258
rect 2365 15206 2377 15258
rect 2429 15206 2441 15258
rect 2493 15206 2505 15258
rect 2557 15206 5951 15258
rect 6003 15206 6015 15258
rect 6067 15206 6079 15258
rect 6131 15206 6143 15258
rect 6195 15206 6207 15258
rect 6259 15206 9653 15258
rect 9705 15206 9717 15258
rect 9769 15206 9781 15258
rect 9833 15206 9845 15258
rect 9897 15206 9909 15258
rect 9961 15206 13355 15258
rect 13407 15206 13419 15258
rect 13471 15206 13483 15258
rect 13535 15206 13547 15258
rect 13599 15206 13611 15258
rect 13663 15206 15364 15258
rect 552 15184 15364 15206
rect 9398 15104 9404 15156
rect 9456 15144 9462 15156
rect 9456 15116 11284 15144
rect 9456 15104 9462 15116
rect 4341 15079 4399 15085
rect 4341 15045 4353 15079
rect 4387 15076 4399 15079
rect 7377 15079 7435 15085
rect 4387 15048 4752 15076
rect 4387 15045 4399 15048
rect 4341 15039 4399 15045
rect 3513 15011 3571 15017
rect 3513 14977 3525 15011
rect 3559 15008 3571 15011
rect 4157 15011 4215 15017
rect 4157 15008 4169 15011
rect 3559 14980 4169 15008
rect 3559 14977 3571 14980
rect 3513 14971 3571 14977
rect 4157 14977 4169 14980
rect 4203 15008 4215 15011
rect 4203 14980 4568 15008
rect 4203 14977 4215 14980
rect 4157 14971 4215 14977
rect 1210 14900 1216 14952
rect 1268 14940 1274 14952
rect 1305 14943 1363 14949
rect 1305 14940 1317 14943
rect 1268 14912 1317 14940
rect 1268 14900 1274 14912
rect 1305 14909 1317 14912
rect 1351 14909 1363 14943
rect 1305 14903 1363 14909
rect 3142 14900 3148 14952
rect 3200 14940 3206 14952
rect 3329 14943 3387 14949
rect 3329 14940 3341 14943
rect 3200 14912 3341 14940
rect 3200 14900 3206 14912
rect 3329 14909 3341 14912
rect 3375 14909 3387 14943
rect 3329 14903 3387 14909
rect 4433 14943 4491 14949
rect 4433 14909 4445 14943
rect 4479 14909 4491 14943
rect 4433 14903 4491 14909
rect 4448 14872 4476 14903
rect 4540 14884 4568 14980
rect 4264 14844 4476 14872
rect 1486 14764 1492 14816
rect 1544 14764 1550 14816
rect 3970 14764 3976 14816
rect 4028 14804 4034 14816
rect 4264 14804 4292 14844
rect 4522 14832 4528 14884
rect 4580 14832 4586 14884
rect 4724 14816 4752 15048
rect 7377 15045 7389 15079
rect 7423 15076 7435 15079
rect 7423 15048 11192 15076
rect 7423 15045 7435 15048
rect 7377 15039 7435 15045
rect 10962 14968 10968 15020
rect 11020 14968 11026 15020
rect 5074 14900 5080 14952
rect 5132 14940 5138 14952
rect 5169 14943 5227 14949
rect 5169 14940 5181 14943
rect 5132 14912 5181 14940
rect 5132 14900 5138 14912
rect 5169 14909 5181 14912
rect 5215 14909 5227 14943
rect 5169 14903 5227 14909
rect 6365 14943 6423 14949
rect 6365 14909 6377 14943
rect 6411 14940 6423 14943
rect 6457 14943 6515 14949
rect 6457 14940 6469 14943
rect 6411 14912 6469 14940
rect 6411 14909 6423 14912
rect 6365 14903 6423 14909
rect 6457 14909 6469 14912
rect 6503 14909 6515 14943
rect 6457 14903 6515 14909
rect 6546 14900 6552 14952
rect 6604 14940 6610 14952
rect 7009 14943 7067 14949
rect 7009 14940 7021 14943
rect 6604 14912 7021 14940
rect 6604 14900 6610 14912
rect 7009 14909 7021 14912
rect 7055 14909 7067 14943
rect 7009 14903 7067 14909
rect 7098 14900 7104 14952
rect 7156 14940 7162 14952
rect 7193 14943 7251 14949
rect 7193 14940 7205 14943
rect 7156 14912 7205 14940
rect 7156 14900 7162 14912
rect 7193 14909 7205 14912
rect 7239 14909 7251 14943
rect 7193 14903 7251 14909
rect 8573 14943 8631 14949
rect 8573 14909 8585 14943
rect 8619 14940 8631 14943
rect 8754 14940 8760 14952
rect 8619 14912 8760 14940
rect 8619 14909 8631 14912
rect 8573 14903 8631 14909
rect 8754 14900 8760 14912
rect 8812 14900 8818 14952
rect 8849 14943 8907 14949
rect 8849 14909 8861 14943
rect 8895 14909 8907 14943
rect 8849 14903 8907 14909
rect 9217 14943 9275 14949
rect 9217 14909 9229 14943
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 5626 14832 5632 14884
rect 5684 14872 5690 14884
rect 8864 14872 8892 14903
rect 5684 14844 8892 14872
rect 9232 14872 9260 14903
rect 9674 14900 9680 14952
rect 9732 14900 9738 14952
rect 11164 14872 11192 15048
rect 11256 14949 11284 15116
rect 11241 14943 11299 14949
rect 11241 14909 11253 14943
rect 11287 14940 11299 14943
rect 12434 14940 12440 14952
rect 11287 14912 12440 14940
rect 11287 14909 11299 14912
rect 11241 14903 11299 14909
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 12802 14900 12808 14952
rect 12860 14940 12866 14952
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 12860 14912 12909 14940
rect 12860 14900 12866 14912
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 11974 14872 11980 14884
rect 9232 14844 10456 14872
rect 11164 14844 11980 14872
rect 5684 14832 5690 14844
rect 10428 14816 10456 14844
rect 11974 14832 11980 14844
rect 12032 14832 12038 14884
rect 4028 14776 4292 14804
rect 4028 14764 4034 14776
rect 4430 14764 4436 14816
rect 4488 14764 4494 14816
rect 4706 14764 4712 14816
rect 4764 14804 4770 14816
rect 5353 14807 5411 14813
rect 5353 14804 5365 14807
rect 4764 14776 5365 14804
rect 4764 14764 4770 14776
rect 5353 14773 5365 14776
rect 5399 14773 5411 14807
rect 5353 14767 5411 14773
rect 6270 14764 6276 14816
rect 6328 14764 6334 14816
rect 8754 14764 8760 14816
rect 8812 14764 8818 14816
rect 9033 14807 9091 14813
rect 9033 14773 9045 14807
rect 9079 14804 9091 14807
rect 9306 14804 9312 14816
rect 9079 14776 9312 14804
rect 9079 14773 9091 14776
rect 9033 14767 9091 14773
rect 9306 14764 9312 14776
rect 9364 14764 9370 14816
rect 10318 14764 10324 14816
rect 10376 14764 10382 14816
rect 10410 14764 10416 14816
rect 10468 14764 10474 14816
rect 11882 14764 11888 14816
rect 11940 14764 11946 14816
rect 13078 14764 13084 14816
rect 13136 14764 13142 14816
rect 552 14714 15520 14736
rect 552 14662 4100 14714
rect 4152 14662 4164 14714
rect 4216 14662 4228 14714
rect 4280 14662 4292 14714
rect 4344 14662 4356 14714
rect 4408 14662 7802 14714
rect 7854 14662 7866 14714
rect 7918 14662 7930 14714
rect 7982 14662 7994 14714
rect 8046 14662 8058 14714
rect 8110 14662 11504 14714
rect 11556 14662 11568 14714
rect 11620 14662 11632 14714
rect 11684 14662 11696 14714
rect 11748 14662 11760 14714
rect 11812 14662 15206 14714
rect 15258 14662 15270 14714
rect 15322 14662 15334 14714
rect 15386 14662 15398 14714
rect 15450 14662 15462 14714
rect 15514 14662 15520 14714
rect 552 14640 15520 14662
rect 1486 14560 1492 14612
rect 1544 14560 1550 14612
rect 3970 14560 3976 14612
rect 4028 14600 4034 14612
rect 4801 14603 4859 14609
rect 4028 14572 4108 14600
rect 4028 14560 4034 14572
rect 1504 14464 1532 14560
rect 3697 14467 3755 14473
rect 3697 14464 3709 14467
rect 1504 14436 3709 14464
rect 3697 14433 3709 14436
rect 3743 14433 3755 14467
rect 3697 14427 3755 14433
rect 3605 14399 3663 14405
rect 3605 14365 3617 14399
rect 3651 14365 3663 14399
rect 3605 14359 3663 14365
rect 3620 14260 3648 14359
rect 3712 14328 3740 14427
rect 4080 14405 4108 14572
rect 4801 14569 4813 14603
rect 4847 14600 4859 14603
rect 8662 14600 8668 14612
rect 4847 14572 8668 14600
rect 4847 14569 4859 14572
rect 4801 14563 4859 14569
rect 8662 14560 8668 14572
rect 8720 14560 8726 14612
rect 8754 14560 8760 14612
rect 8812 14600 8818 14612
rect 9493 14603 9551 14609
rect 9493 14600 9505 14603
rect 8812 14572 9505 14600
rect 8812 14560 8818 14572
rect 9493 14569 9505 14572
rect 9539 14569 9551 14603
rect 9493 14563 9551 14569
rect 9585 14603 9643 14609
rect 9585 14569 9597 14603
rect 9631 14600 9643 14603
rect 9674 14600 9680 14612
rect 9631 14572 9680 14600
rect 9631 14569 9643 14572
rect 9585 14563 9643 14569
rect 4522 14532 4528 14544
rect 4356 14504 4528 14532
rect 4356 14473 4384 14504
rect 4522 14492 4528 14504
rect 4580 14532 4586 14544
rect 5261 14535 5319 14541
rect 4580 14504 5212 14532
rect 4580 14492 4586 14504
rect 4157 14467 4215 14473
rect 4157 14433 4169 14467
rect 4203 14433 4215 14467
rect 4157 14427 4215 14433
rect 4341 14467 4399 14473
rect 4341 14433 4353 14467
rect 4387 14433 4399 14467
rect 4341 14427 4399 14433
rect 4065 14399 4123 14405
rect 4065 14365 4077 14399
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 4172 14396 4200 14427
rect 4430 14424 4436 14476
rect 4488 14424 4494 14476
rect 4614 14424 4620 14476
rect 4672 14424 4678 14476
rect 5077 14467 5135 14473
rect 5077 14464 5089 14467
rect 5000 14436 5089 14464
rect 4172 14368 4660 14396
rect 4172 14328 4200 14368
rect 3712 14300 4200 14328
rect 4522 14288 4528 14340
rect 4580 14288 4586 14340
rect 4632 14328 4660 14368
rect 5000 14328 5028 14436
rect 5077 14433 5089 14436
rect 5123 14433 5135 14467
rect 5184 14464 5212 14504
rect 5261 14501 5273 14535
rect 5307 14532 5319 14535
rect 5813 14535 5871 14541
rect 5813 14532 5825 14535
rect 5307 14504 5825 14532
rect 5307 14501 5319 14504
rect 5261 14495 5319 14501
rect 5813 14501 5825 14504
rect 5859 14501 5871 14535
rect 5813 14495 5871 14501
rect 7116 14504 7696 14532
rect 7116 14476 7144 14504
rect 5350 14464 5356 14476
rect 5184 14436 5356 14464
rect 5077 14427 5135 14433
rect 5350 14424 5356 14436
rect 5408 14424 5414 14476
rect 5442 14424 5448 14476
rect 5500 14424 5506 14476
rect 6089 14467 6147 14473
rect 6089 14433 6101 14467
rect 6135 14433 6147 14467
rect 6089 14427 6147 14433
rect 5813 14399 5871 14405
rect 5813 14396 5825 14399
rect 5736 14368 5825 14396
rect 5166 14328 5172 14340
rect 4632 14300 5172 14328
rect 5166 14288 5172 14300
rect 5224 14288 5230 14340
rect 5626 14288 5632 14340
rect 5684 14288 5690 14340
rect 5736 14328 5764 14368
rect 5813 14365 5825 14368
rect 5859 14365 5871 14399
rect 6104 14396 6132 14427
rect 7098 14424 7104 14476
rect 7156 14424 7162 14476
rect 7397 14467 7455 14473
rect 7397 14433 7409 14467
rect 7443 14464 7455 14467
rect 7558 14464 7564 14476
rect 7443 14436 7564 14464
rect 7443 14433 7455 14436
rect 7397 14427 7455 14433
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 7668 14473 7696 14504
rect 9398 14492 9404 14544
rect 9456 14492 9462 14544
rect 7653 14467 7711 14473
rect 7653 14433 7665 14467
rect 7699 14464 7711 14467
rect 7745 14467 7803 14473
rect 7745 14464 7757 14467
rect 7699 14436 7757 14464
rect 7699 14433 7711 14436
rect 7653 14427 7711 14433
rect 7745 14433 7757 14436
rect 7791 14433 7803 14467
rect 7745 14427 7803 14433
rect 8012 14467 8070 14473
rect 8012 14433 8024 14467
rect 8058 14464 8070 14467
rect 8386 14464 8392 14476
rect 8058 14436 8392 14464
rect 8058 14433 8070 14436
rect 8012 14427 8070 14433
rect 8386 14424 8392 14436
rect 8444 14424 8450 14476
rect 6362 14396 6368 14408
rect 6104 14368 6368 14396
rect 5813 14359 5871 14365
rect 6362 14356 6368 14368
rect 6420 14356 6426 14408
rect 9416 14405 9444 14492
rect 9401 14399 9459 14405
rect 9401 14365 9413 14399
rect 9447 14365 9459 14399
rect 9401 14359 9459 14365
rect 6273 14331 6331 14337
rect 6273 14328 6285 14331
rect 5736 14300 6285 14328
rect 5736 14260 5764 14300
rect 6273 14297 6285 14300
rect 6319 14328 6331 14331
rect 6546 14328 6552 14340
rect 6319 14300 6552 14328
rect 6319 14297 6331 14300
rect 6273 14291 6331 14297
rect 6546 14288 6552 14300
rect 6604 14288 6610 14340
rect 9125 14331 9183 14337
rect 9125 14297 9137 14331
rect 9171 14328 9183 14331
rect 9600 14328 9628 14563
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 10318 14560 10324 14612
rect 10376 14560 10382 14612
rect 13814 14600 13820 14612
rect 11992 14572 13820 14600
rect 10229 14467 10287 14473
rect 10229 14433 10241 14467
rect 10275 14464 10287 14467
rect 10336 14464 10364 14560
rect 11992 14532 12020 14572
rect 13814 14560 13820 14572
rect 13872 14560 13878 14612
rect 14093 14535 14151 14541
rect 14093 14532 14105 14535
rect 10275 14436 10364 14464
rect 11164 14504 12020 14532
rect 12926 14504 14105 14532
rect 10275 14433 10287 14436
rect 10229 14427 10287 14433
rect 9171 14300 9628 14328
rect 9953 14331 10011 14337
rect 9171 14297 9183 14300
rect 9125 14291 9183 14297
rect 9953 14297 9965 14331
rect 9999 14328 10011 14331
rect 11164 14328 11192 14504
rect 14093 14501 14105 14504
rect 14139 14501 14151 14535
rect 14093 14495 14151 14501
rect 11425 14467 11483 14473
rect 11425 14464 11437 14467
rect 11348 14436 11437 14464
rect 11348 14408 11376 14436
rect 11425 14433 11437 14436
rect 11471 14433 11483 14467
rect 11425 14427 11483 14433
rect 13078 14424 13084 14476
rect 13136 14464 13142 14476
rect 14001 14467 14059 14473
rect 14001 14464 14013 14467
rect 13136 14436 14013 14464
rect 13136 14424 13142 14436
rect 14001 14433 14013 14436
rect 14047 14433 14059 14467
rect 14001 14427 14059 14433
rect 11330 14356 11336 14408
rect 11388 14356 11394 14408
rect 11701 14399 11759 14405
rect 11701 14365 11713 14399
rect 11747 14396 11759 14399
rect 11790 14396 11796 14408
rect 11747 14368 11796 14396
rect 11747 14365 11759 14368
rect 11701 14359 11759 14365
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 13173 14399 13231 14405
rect 13173 14365 13185 14399
rect 13219 14396 13231 14399
rect 13817 14399 13875 14405
rect 13817 14396 13829 14399
rect 13219 14368 13829 14396
rect 13219 14365 13231 14368
rect 13173 14359 13231 14365
rect 13817 14365 13829 14368
rect 13863 14365 13875 14399
rect 13817 14359 13875 14365
rect 9999 14300 11192 14328
rect 9999 14297 10011 14300
rect 9953 14291 10011 14297
rect 3620 14232 5764 14260
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 5997 14263 6055 14269
rect 5997 14260 6009 14263
rect 5868 14232 6009 14260
rect 5868 14220 5874 14232
rect 5997 14229 6009 14232
rect 6043 14229 6055 14263
rect 5997 14223 6055 14229
rect 7374 14220 7380 14272
rect 7432 14260 7438 14272
rect 9306 14260 9312 14272
rect 7432 14232 9312 14260
rect 7432 14220 7438 14232
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 9490 14220 9496 14272
rect 9548 14260 9554 14272
rect 10137 14263 10195 14269
rect 10137 14260 10149 14263
rect 9548 14232 10149 14260
rect 9548 14220 9554 14232
rect 10137 14229 10149 14232
rect 10183 14229 10195 14263
rect 10137 14223 10195 14229
rect 10410 14220 10416 14272
rect 10468 14260 10474 14272
rect 13188 14260 13216 14359
rect 10468 14232 13216 14260
rect 10468 14220 10474 14232
rect 13262 14220 13268 14272
rect 13320 14220 13326 14272
rect 552 14170 15364 14192
rect 552 14118 2249 14170
rect 2301 14118 2313 14170
rect 2365 14118 2377 14170
rect 2429 14118 2441 14170
rect 2493 14118 2505 14170
rect 2557 14118 5951 14170
rect 6003 14118 6015 14170
rect 6067 14118 6079 14170
rect 6131 14118 6143 14170
rect 6195 14118 6207 14170
rect 6259 14118 9653 14170
rect 9705 14118 9717 14170
rect 9769 14118 9781 14170
rect 9833 14118 9845 14170
rect 9897 14118 9909 14170
rect 9961 14118 13355 14170
rect 13407 14118 13419 14170
rect 13471 14118 13483 14170
rect 13535 14118 13547 14170
rect 13599 14118 13611 14170
rect 13663 14118 15364 14170
rect 552 14096 15364 14118
rect 3970 14016 3976 14068
rect 4028 14016 4034 14068
rect 4522 14016 4528 14068
rect 4580 14056 4586 14068
rect 4709 14059 4767 14065
rect 4709 14056 4721 14059
rect 4580 14028 4721 14056
rect 4580 14016 4586 14028
rect 4709 14025 4721 14028
rect 4755 14025 4767 14059
rect 4709 14019 4767 14025
rect 5442 14016 5448 14068
rect 5500 14056 5506 14068
rect 5629 14059 5687 14065
rect 5629 14056 5641 14059
rect 5500 14028 5641 14056
rect 5500 14016 5506 14028
rect 5629 14025 5641 14028
rect 5675 14025 5687 14059
rect 5629 14019 5687 14025
rect 6270 14016 6276 14068
rect 6328 14016 6334 14068
rect 7190 14056 7196 14068
rect 6564 14028 7196 14056
rect 3988 13920 4016 14016
rect 4341 13991 4399 13997
rect 4341 13957 4353 13991
rect 4387 13988 4399 13991
rect 4387 13960 4752 13988
rect 4387 13957 4399 13960
rect 4341 13951 4399 13957
rect 3988 13892 4568 13920
rect 4540 13861 4568 13892
rect 4724 13864 4752 13960
rect 5166 13880 5172 13932
rect 5224 13920 5230 13932
rect 6288 13929 6316 14016
rect 6181 13923 6239 13929
rect 6181 13920 6193 13923
rect 5224 13892 6193 13920
rect 5224 13880 5230 13892
rect 6181 13889 6193 13892
rect 6227 13889 6239 13923
rect 6181 13883 6239 13889
rect 6273 13923 6331 13929
rect 6273 13889 6285 13923
rect 6319 13920 6331 13923
rect 6319 13892 6500 13920
rect 6319 13889 6331 13892
rect 6273 13883 6331 13889
rect 4249 13855 4307 13861
rect 4249 13821 4261 13855
rect 4295 13821 4307 13855
rect 4249 13815 4307 13821
rect 4525 13855 4583 13861
rect 4525 13821 4537 13855
rect 4571 13821 4583 13855
rect 4525 13815 4583 13821
rect 4264 13784 4292 13815
rect 4706 13812 4712 13864
rect 4764 13812 4770 13864
rect 5258 13812 5264 13864
rect 5316 13812 5322 13864
rect 5810 13855 5868 13861
rect 5810 13821 5822 13855
rect 5856 13852 5868 13855
rect 6362 13852 6368 13864
rect 5856 13824 6368 13852
rect 5856 13821 5868 13824
rect 5810 13815 5868 13821
rect 5276 13784 5304 13812
rect 4264 13756 5304 13784
rect 5350 13676 5356 13728
rect 5408 13716 5414 13728
rect 5810 13716 5816 13728
rect 5408 13688 5816 13716
rect 5408 13676 5414 13688
rect 5810 13676 5816 13688
rect 5868 13676 5874 13728
rect 6288 13716 6316 13824
rect 6362 13812 6368 13824
rect 6420 13812 6426 13864
rect 6472 13784 6500 13892
rect 6564 13861 6592 14028
rect 7190 14016 7196 14028
rect 7248 14056 7254 14068
rect 7248 14028 7512 14056
rect 7248 14016 7254 14028
rect 6825 13991 6883 13997
rect 6825 13957 6837 13991
rect 6871 13957 6883 13991
rect 7374 13988 7380 14000
rect 6825 13951 6883 13957
rect 7208 13960 7380 13988
rect 6840 13920 6868 13951
rect 7009 13923 7067 13929
rect 7009 13920 7021 13923
rect 6840 13892 7021 13920
rect 7009 13889 7021 13892
rect 7055 13889 7067 13923
rect 7009 13883 7067 13889
rect 6549 13855 6607 13861
rect 6549 13821 6561 13855
rect 6595 13821 6607 13855
rect 6549 13815 6607 13821
rect 6641 13855 6699 13861
rect 6641 13821 6653 13855
rect 6687 13821 6699 13855
rect 7208 13852 7236 13960
rect 7374 13948 7380 13960
rect 7432 13948 7438 14000
rect 7484 13920 7512 14028
rect 7558 14016 7564 14068
rect 7616 14056 7622 14068
rect 7653 14059 7711 14065
rect 7653 14056 7665 14059
rect 7616 14028 7665 14056
rect 7616 14016 7622 14028
rect 7653 14025 7665 14028
rect 7699 14025 7711 14059
rect 7653 14019 7711 14025
rect 8386 14016 8392 14068
rect 8444 14016 8450 14068
rect 9398 14016 9404 14068
rect 9456 14016 9462 14068
rect 10410 14016 10416 14068
rect 10468 14016 10474 14068
rect 11422 14016 11428 14068
rect 11480 14056 11486 14068
rect 11885 14059 11943 14065
rect 11885 14056 11897 14059
rect 11480 14028 11897 14056
rect 11480 14016 11486 14028
rect 11885 14025 11897 14028
rect 11931 14025 11943 14059
rect 11885 14019 11943 14025
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 12713 14059 12771 14065
rect 12713 14056 12725 14059
rect 12492 14028 12725 14056
rect 12492 14016 12498 14028
rect 12713 14025 12725 14028
rect 12759 14025 12771 14059
rect 12713 14019 12771 14025
rect 9416 13988 9444 14016
rect 9416 13960 9628 13988
rect 7837 13923 7895 13929
rect 7837 13920 7849 13923
rect 7484 13892 7849 13920
rect 7837 13889 7849 13892
rect 7883 13889 7895 13923
rect 9125 13923 9183 13929
rect 9125 13920 9137 13923
rect 7837 13883 7895 13889
rect 8588 13892 9137 13920
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 6641 13815 6699 13821
rect 6840 13824 7236 13852
rect 7392 13824 7757 13852
rect 6656 13784 6684 13815
rect 6840 13793 6868 13824
rect 6472 13756 6684 13784
rect 6825 13787 6883 13793
rect 6825 13753 6837 13787
rect 6871 13753 6883 13787
rect 6825 13747 6883 13753
rect 6730 13716 6736 13728
rect 6288 13688 6736 13716
rect 6730 13676 6736 13688
rect 6788 13716 6794 13728
rect 7392 13716 7420 13824
rect 7745 13821 7757 13824
rect 7791 13821 7803 13855
rect 7745 13815 7803 13821
rect 7929 13855 7987 13861
rect 7929 13821 7941 13855
rect 7975 13852 7987 13855
rect 8202 13852 8208 13864
rect 7975 13824 8208 13852
rect 7975 13821 7987 13824
rect 7929 13815 7987 13821
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 8588 13861 8616 13892
rect 9125 13889 9137 13892
rect 9171 13889 9183 13923
rect 9490 13920 9496 13932
rect 9125 13883 9183 13889
rect 9232 13892 9496 13920
rect 8573 13855 8631 13861
rect 8573 13821 8585 13855
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 8662 13812 8668 13864
rect 8720 13852 8726 13864
rect 8849 13855 8907 13861
rect 8849 13852 8861 13855
rect 8720 13824 8861 13852
rect 8720 13812 8726 13824
rect 8849 13821 8861 13824
rect 8895 13852 8907 13855
rect 9033 13855 9091 13861
rect 8895 13824 8984 13852
rect 8895 13821 8907 13824
rect 8849 13815 8907 13821
rect 8956 13784 8984 13824
rect 9033 13821 9045 13855
rect 9079 13852 9091 13855
rect 9232 13852 9260 13892
rect 9416 13861 9444 13892
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 9600 13861 9628 13960
rect 9079 13824 9260 13852
rect 9309 13855 9367 13861
rect 9079 13821 9091 13824
rect 9033 13815 9091 13821
rect 9309 13821 9321 13855
rect 9355 13821 9367 13855
rect 9309 13815 9367 13821
rect 9401 13855 9459 13861
rect 9401 13821 9413 13855
rect 9447 13821 9459 13855
rect 9401 13815 9459 13821
rect 9585 13855 9643 13861
rect 9585 13821 9597 13855
rect 9631 13821 9643 13855
rect 9585 13815 9643 13821
rect 9677 13855 9735 13861
rect 9677 13821 9689 13855
rect 9723 13852 9735 13855
rect 10428 13852 10456 14016
rect 14734 13988 14740 14000
rect 11808 13960 14740 13988
rect 11808 13861 11836 13960
rect 14734 13948 14740 13960
rect 14792 13948 14798 14000
rect 11974 13880 11980 13932
rect 12032 13920 12038 13932
rect 12345 13923 12403 13929
rect 12345 13920 12357 13923
rect 12032 13892 12357 13920
rect 12032 13880 12038 13892
rect 12345 13889 12357 13892
rect 12391 13889 12403 13923
rect 12345 13883 12403 13889
rect 12434 13880 12440 13932
rect 12492 13880 12498 13932
rect 13262 13920 13268 13932
rect 13004 13892 13268 13920
rect 9723 13824 10456 13852
rect 11793 13855 11851 13861
rect 9723 13821 9735 13824
rect 9677 13815 9735 13821
rect 11793 13821 11805 13855
rect 11839 13821 11851 13855
rect 11793 13815 11851 13821
rect 9324 13784 9352 13815
rect 11882 13812 11888 13864
rect 11940 13852 11946 13864
rect 13004 13861 13032 13892
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 12713 13855 12771 13861
rect 12713 13852 12725 13855
rect 11940 13824 12725 13852
rect 11940 13812 11946 13824
rect 12713 13821 12725 13824
rect 12759 13821 12771 13855
rect 12713 13815 12771 13821
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 12989 13855 13047 13861
rect 12989 13821 13001 13855
rect 13035 13821 13047 13855
rect 13725 13855 13783 13861
rect 13725 13852 13737 13855
rect 12989 13815 13047 13821
rect 13188 13824 13737 13852
rect 9766 13784 9772 13796
rect 8956 13756 9772 13784
rect 9766 13744 9772 13756
rect 9824 13744 9830 13796
rect 11238 13744 11244 13796
rect 11296 13784 11302 13796
rect 12912 13784 12940 13815
rect 11296 13756 12940 13784
rect 11296 13744 11302 13756
rect 6788 13688 7420 13716
rect 6788 13676 6794 13688
rect 10042 13676 10048 13728
rect 10100 13716 10106 13728
rect 10321 13719 10379 13725
rect 10321 13716 10333 13719
rect 10100 13688 10333 13716
rect 10100 13676 10106 13688
rect 10321 13685 10333 13688
rect 10367 13685 10379 13719
rect 10321 13679 10379 13685
rect 12250 13676 12256 13728
rect 12308 13676 12314 13728
rect 13188 13725 13216 13824
rect 13725 13821 13737 13824
rect 13771 13821 13783 13855
rect 13725 13815 13783 13821
rect 13173 13719 13231 13725
rect 13173 13685 13185 13719
rect 13219 13685 13231 13719
rect 13173 13679 13231 13685
rect 13262 13676 13268 13728
rect 13320 13716 13326 13728
rect 13541 13719 13599 13725
rect 13541 13716 13553 13719
rect 13320 13688 13553 13716
rect 13320 13676 13326 13688
rect 13541 13685 13553 13688
rect 13587 13685 13599 13719
rect 13541 13679 13599 13685
rect 552 13626 15520 13648
rect 552 13574 4100 13626
rect 4152 13574 4164 13626
rect 4216 13574 4228 13626
rect 4280 13574 4292 13626
rect 4344 13574 4356 13626
rect 4408 13574 7802 13626
rect 7854 13574 7866 13626
rect 7918 13574 7930 13626
rect 7982 13574 7994 13626
rect 8046 13574 8058 13626
rect 8110 13574 11504 13626
rect 11556 13574 11568 13626
rect 11620 13574 11632 13626
rect 11684 13574 11696 13626
rect 11748 13574 11760 13626
rect 11812 13574 15206 13626
rect 15258 13574 15270 13626
rect 15322 13574 15334 13626
rect 15386 13574 15398 13626
rect 15450 13574 15462 13626
rect 15514 13574 15520 13626
rect 552 13552 15520 13574
rect 4614 13472 4620 13524
rect 4672 13512 4678 13524
rect 4709 13515 4767 13521
rect 4709 13512 4721 13515
rect 4672 13484 4721 13512
rect 4672 13472 4678 13484
rect 4709 13481 4721 13484
rect 4755 13481 4767 13515
rect 4709 13475 4767 13481
rect 10321 13515 10379 13521
rect 10321 13481 10333 13515
rect 10367 13512 10379 13515
rect 11238 13512 11244 13524
rect 10367 13484 11244 13512
rect 10367 13481 10379 13484
rect 10321 13475 10379 13481
rect 11238 13472 11244 13484
rect 11296 13472 11302 13524
rect 12250 13472 12256 13524
rect 12308 13472 12314 13524
rect 7561 13447 7619 13453
rect 7561 13413 7573 13447
rect 7607 13444 7619 13447
rect 10042 13444 10048 13456
rect 7607 13416 10048 13444
rect 7607 13413 7619 13416
rect 7561 13407 7619 13413
rect 10042 13404 10048 13416
rect 10100 13444 10106 13456
rect 10965 13447 11023 13453
rect 10965 13444 10977 13447
rect 10100 13416 10977 13444
rect 10100 13404 10106 13416
rect 10965 13413 10977 13416
rect 11011 13413 11023 13447
rect 10965 13407 11023 13413
rect 5077 13379 5135 13385
rect 5077 13345 5089 13379
rect 5123 13376 5135 13379
rect 5350 13376 5356 13388
rect 5123 13348 5356 13376
rect 5123 13345 5135 13348
rect 5077 13339 5135 13345
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 7374 13336 7380 13388
rect 7432 13376 7438 13388
rect 7653 13379 7711 13385
rect 7653 13376 7665 13379
rect 7432 13348 7665 13376
rect 7432 13336 7438 13348
rect 7653 13345 7665 13348
rect 7699 13345 7711 13379
rect 7653 13339 7711 13345
rect 9766 13336 9772 13388
rect 9824 13376 9830 13388
rect 10137 13379 10195 13385
rect 10137 13376 10149 13379
rect 9824 13348 10149 13376
rect 9824 13336 9830 13348
rect 10137 13345 10149 13348
rect 10183 13376 10195 13379
rect 10413 13379 10471 13385
rect 10413 13376 10425 13379
rect 10183 13348 10425 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 10413 13345 10425 13348
rect 10459 13345 10471 13379
rect 10413 13339 10471 13345
rect 10597 13379 10655 13385
rect 10597 13345 10609 13379
rect 10643 13376 10655 13379
rect 10870 13376 10876 13388
rect 10643 13348 10876 13376
rect 10643 13345 10655 13348
rect 10597 13339 10655 13345
rect 10870 13336 10876 13348
rect 10928 13376 10934 13388
rect 12268 13376 12296 13472
rect 10928 13348 12296 13376
rect 10928 13336 10934 13348
rect 5166 13268 5172 13320
rect 5224 13268 5230 13320
rect 5261 13311 5319 13317
rect 5261 13277 5273 13311
rect 5307 13277 5319 13311
rect 5261 13271 5319 13277
rect 9953 13311 10011 13317
rect 9953 13277 9965 13311
rect 9999 13277 10011 13311
rect 9953 13271 10011 13277
rect 10505 13311 10563 13317
rect 10505 13277 10517 13311
rect 10551 13308 10563 13311
rect 11882 13308 11888 13320
rect 10551 13280 11888 13308
rect 10551 13277 10563 13280
rect 10505 13271 10563 13277
rect 4798 13200 4804 13252
rect 4856 13240 4862 13252
rect 5276 13240 5304 13271
rect 4856 13212 5304 13240
rect 9968 13240 9996 13271
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 10870 13240 10876 13252
rect 9968 13212 10876 13240
rect 4856 13200 4862 13212
rect 10870 13200 10876 13212
rect 10928 13200 10934 13252
rect 6273 13175 6331 13181
rect 6273 13141 6285 13175
rect 6319 13172 6331 13175
rect 7098 13172 7104 13184
rect 6319 13144 7104 13172
rect 6319 13141 6331 13144
rect 6273 13135 6331 13141
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 7834 13132 7840 13184
rect 7892 13132 7898 13184
rect 12250 13132 12256 13184
rect 12308 13132 12314 13184
rect 552 13082 15364 13104
rect 552 13030 2249 13082
rect 2301 13030 2313 13082
rect 2365 13030 2377 13082
rect 2429 13030 2441 13082
rect 2493 13030 2505 13082
rect 2557 13030 5951 13082
rect 6003 13030 6015 13082
rect 6067 13030 6079 13082
rect 6131 13030 6143 13082
rect 6195 13030 6207 13082
rect 6259 13030 9653 13082
rect 9705 13030 9717 13082
rect 9769 13030 9781 13082
rect 9833 13030 9845 13082
rect 9897 13030 9909 13082
rect 9961 13030 13355 13082
rect 13407 13030 13419 13082
rect 13471 13030 13483 13082
rect 13535 13030 13547 13082
rect 13599 13030 13611 13082
rect 13663 13030 15364 13082
rect 552 13008 15364 13030
rect 4706 12928 4712 12980
rect 4764 12928 4770 12980
rect 4798 12928 4804 12980
rect 4856 12928 4862 12980
rect 5166 12928 5172 12980
rect 5224 12968 5230 12980
rect 5445 12971 5503 12977
rect 5445 12968 5457 12971
rect 5224 12940 5457 12968
rect 5224 12928 5230 12940
rect 5445 12937 5457 12940
rect 5491 12937 5503 12971
rect 5445 12931 5503 12937
rect 5629 12971 5687 12977
rect 5629 12937 5641 12971
rect 5675 12937 5687 12971
rect 5629 12931 5687 12937
rect 4724 12900 4752 12928
rect 5644 12900 5672 12931
rect 6730 12928 6736 12980
rect 6788 12928 6794 12980
rect 10870 12928 10876 12980
rect 10928 12968 10934 12980
rect 10965 12971 11023 12977
rect 10965 12968 10977 12971
rect 10928 12940 10977 12968
rect 10928 12928 10934 12940
rect 10965 12937 10977 12940
rect 11011 12937 11023 12971
rect 10965 12931 11023 12937
rect 4724 12872 5672 12900
rect 5077 12835 5135 12841
rect 5077 12801 5089 12835
rect 5123 12801 5135 12835
rect 5077 12795 5135 12801
rect 5092 12696 5120 12795
rect 7098 12792 7104 12844
rect 7156 12792 7162 12844
rect 5169 12767 5227 12773
rect 5169 12733 5181 12767
rect 5215 12764 5227 12767
rect 5258 12764 5264 12776
rect 5215 12736 5264 12764
rect 5215 12733 5227 12736
rect 5169 12727 5227 12733
rect 5258 12724 5264 12736
rect 5316 12724 5322 12776
rect 5902 12724 5908 12776
rect 5960 12764 5966 12776
rect 6641 12767 6699 12773
rect 5960 12736 6500 12764
rect 5960 12724 5966 12736
rect 6472 12705 6500 12736
rect 6641 12733 6653 12767
rect 6687 12764 6699 12767
rect 7006 12764 7012 12776
rect 6687 12736 7012 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 7116 12764 7144 12792
rect 8113 12767 8171 12773
rect 8113 12764 8125 12767
rect 7116 12736 8125 12764
rect 8113 12733 8125 12736
rect 8159 12733 8171 12767
rect 8113 12727 8171 12733
rect 9769 12767 9827 12773
rect 9769 12733 9781 12767
rect 9815 12764 9827 12767
rect 11330 12764 11336 12776
rect 9815 12736 11336 12764
rect 9815 12733 9827 12736
rect 9769 12727 9827 12733
rect 11330 12724 11336 12736
rect 11388 12764 11394 12776
rect 12250 12764 12256 12776
rect 11388 12736 12256 12764
rect 11388 12724 11394 12736
rect 12250 12724 12256 12736
rect 12308 12764 12314 12776
rect 12345 12767 12403 12773
rect 12345 12764 12357 12767
rect 12308 12736 12357 12764
rect 12308 12724 12314 12736
rect 12345 12733 12357 12736
rect 12391 12733 12403 12767
rect 12345 12727 12403 12733
rect 6273 12699 6331 12705
rect 6273 12696 6285 12699
rect 5092 12668 6285 12696
rect 6273 12665 6285 12668
rect 6319 12665 6331 12699
rect 6273 12659 6331 12665
rect 6457 12699 6515 12705
rect 6457 12665 6469 12699
rect 6503 12696 6515 12699
rect 6503 12668 7052 12696
rect 6503 12665 6515 12668
rect 6457 12659 6515 12665
rect 6288 12628 6316 12659
rect 6730 12628 6736 12640
rect 6288 12600 6736 12628
rect 6730 12588 6736 12600
rect 6788 12588 6794 12640
rect 7024 12628 7052 12668
rect 7834 12656 7840 12708
rect 7892 12705 7898 12708
rect 7892 12696 7904 12705
rect 7892 12668 7937 12696
rect 7892 12659 7904 12668
rect 7892 12656 7898 12659
rect 9398 12656 9404 12708
rect 9456 12696 9462 12708
rect 9502 12699 9560 12705
rect 9502 12696 9514 12699
rect 9456 12668 9514 12696
rect 9456 12656 9462 12668
rect 9502 12665 9514 12668
rect 9548 12665 9560 12699
rect 9502 12659 9560 12665
rect 12100 12699 12158 12705
rect 12100 12665 12112 12699
rect 12146 12696 12158 12699
rect 13262 12696 13268 12708
rect 12146 12668 13268 12696
rect 12146 12665 12158 12668
rect 12100 12659 12158 12665
rect 13262 12656 13268 12668
rect 13320 12656 13326 12708
rect 8386 12628 8392 12640
rect 7024 12600 8392 12628
rect 8386 12588 8392 12600
rect 8444 12588 8450 12640
rect 552 12538 15520 12560
rect 552 12486 4100 12538
rect 4152 12486 4164 12538
rect 4216 12486 4228 12538
rect 4280 12486 4292 12538
rect 4344 12486 4356 12538
rect 4408 12486 7802 12538
rect 7854 12486 7866 12538
rect 7918 12486 7930 12538
rect 7982 12486 7994 12538
rect 8046 12486 8058 12538
rect 8110 12486 11504 12538
rect 11556 12486 11568 12538
rect 11620 12486 11632 12538
rect 11684 12486 11696 12538
rect 11748 12486 11760 12538
rect 11812 12486 15206 12538
rect 15258 12486 15270 12538
rect 15322 12486 15334 12538
rect 15386 12486 15398 12538
rect 15450 12486 15462 12538
rect 15514 12486 15520 12538
rect 552 12464 15520 12486
rect 4706 12384 4712 12436
rect 4764 12384 4770 12436
rect 5350 12384 5356 12436
rect 5408 12384 5414 12436
rect 7009 12427 7067 12433
rect 7009 12393 7021 12427
rect 7055 12424 7067 12427
rect 7098 12424 7104 12436
rect 7055 12396 7104 12424
rect 7055 12393 7067 12396
rect 7009 12387 7067 12393
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 7190 12384 7196 12436
rect 7248 12384 7254 12436
rect 8202 12384 8208 12436
rect 8260 12424 8266 12436
rect 9125 12427 9183 12433
rect 9125 12424 9137 12427
rect 8260 12396 9137 12424
rect 8260 12384 8266 12396
rect 9125 12393 9137 12396
rect 9171 12393 9183 12427
rect 9125 12387 9183 12393
rect 9309 12427 9367 12433
rect 9309 12393 9321 12427
rect 9355 12424 9367 12427
rect 9398 12424 9404 12436
rect 9355 12396 9404 12424
rect 9355 12393 9367 12396
rect 9309 12387 9367 12393
rect 4724 12288 4752 12384
rect 4893 12291 4951 12297
rect 4893 12288 4905 12291
rect 4724 12260 4905 12288
rect 4893 12257 4905 12260
rect 4939 12257 4951 12291
rect 4893 12251 4951 12257
rect 8386 12248 8392 12300
rect 8444 12288 8450 12300
rect 8481 12291 8539 12297
rect 8481 12288 8493 12291
rect 8444 12260 8493 12288
rect 8444 12248 8450 12260
rect 8481 12257 8493 12260
rect 8527 12257 8539 12291
rect 9140 12288 9168 12387
rect 9398 12384 9404 12396
rect 9456 12384 9462 12436
rect 9217 12291 9275 12297
rect 9217 12288 9229 12291
rect 9140 12260 9229 12288
rect 8481 12251 8539 12257
rect 9217 12257 9229 12260
rect 9263 12257 9275 12291
rect 9217 12251 9275 12257
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 9401 12291 9459 12297
rect 9401 12288 9413 12291
rect 9364 12260 9413 12288
rect 9364 12248 9370 12260
rect 9401 12257 9413 12260
rect 9447 12257 9459 12291
rect 9401 12251 9459 12257
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 14553 12291 14611 12297
rect 14553 12288 14565 12291
rect 13872 12260 14565 12288
rect 13872 12248 13878 12260
rect 14553 12257 14565 12260
rect 14599 12257 14611 12291
rect 14553 12251 14611 12257
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 9324 12220 9352 12248
rect 6687 12192 9352 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 5169 12087 5227 12093
rect 5169 12053 5181 12087
rect 5215 12084 5227 12087
rect 5810 12084 5816 12096
rect 5215 12056 5816 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 7006 12044 7012 12096
rect 7064 12044 7070 12096
rect 14734 12044 14740 12096
rect 14792 12044 14798 12096
rect 552 11994 15364 12016
rect 552 11942 2249 11994
rect 2301 11942 2313 11994
rect 2365 11942 2377 11994
rect 2429 11942 2441 11994
rect 2493 11942 2505 11994
rect 2557 11942 5951 11994
rect 6003 11942 6015 11994
rect 6067 11942 6079 11994
rect 6131 11942 6143 11994
rect 6195 11942 6207 11994
rect 6259 11942 9653 11994
rect 9705 11942 9717 11994
rect 9769 11942 9781 11994
rect 9833 11942 9845 11994
rect 9897 11942 9909 11994
rect 9961 11942 13355 11994
rect 13407 11942 13419 11994
rect 13471 11942 13483 11994
rect 13535 11942 13547 11994
rect 13599 11942 13611 11994
rect 13663 11942 15364 11994
rect 552 11920 15364 11942
rect 552 11450 15520 11472
rect 552 11398 4100 11450
rect 4152 11398 4164 11450
rect 4216 11398 4228 11450
rect 4280 11398 4292 11450
rect 4344 11398 4356 11450
rect 4408 11398 7802 11450
rect 7854 11398 7866 11450
rect 7918 11398 7930 11450
rect 7982 11398 7994 11450
rect 8046 11398 8058 11450
rect 8110 11398 11504 11450
rect 11556 11398 11568 11450
rect 11620 11398 11632 11450
rect 11684 11398 11696 11450
rect 11748 11398 11760 11450
rect 11812 11398 15206 11450
rect 15258 11398 15270 11450
rect 15322 11398 15334 11450
rect 15386 11398 15398 11450
rect 15450 11398 15462 11450
rect 15514 11398 15520 11450
rect 552 11376 15520 11398
rect 552 10906 15364 10928
rect 552 10854 2249 10906
rect 2301 10854 2313 10906
rect 2365 10854 2377 10906
rect 2429 10854 2441 10906
rect 2493 10854 2505 10906
rect 2557 10854 5951 10906
rect 6003 10854 6015 10906
rect 6067 10854 6079 10906
rect 6131 10854 6143 10906
rect 6195 10854 6207 10906
rect 6259 10854 9653 10906
rect 9705 10854 9717 10906
rect 9769 10854 9781 10906
rect 9833 10854 9845 10906
rect 9897 10854 9909 10906
rect 9961 10854 13355 10906
rect 13407 10854 13419 10906
rect 13471 10854 13483 10906
rect 13535 10854 13547 10906
rect 13599 10854 13611 10906
rect 13663 10854 15364 10906
rect 552 10832 15364 10854
rect 552 10362 15520 10384
rect 552 10310 4100 10362
rect 4152 10310 4164 10362
rect 4216 10310 4228 10362
rect 4280 10310 4292 10362
rect 4344 10310 4356 10362
rect 4408 10310 7802 10362
rect 7854 10310 7866 10362
rect 7918 10310 7930 10362
rect 7982 10310 7994 10362
rect 8046 10310 8058 10362
rect 8110 10310 11504 10362
rect 11556 10310 11568 10362
rect 11620 10310 11632 10362
rect 11684 10310 11696 10362
rect 11748 10310 11760 10362
rect 11812 10310 15206 10362
rect 15258 10310 15270 10362
rect 15322 10310 15334 10362
rect 15386 10310 15398 10362
rect 15450 10310 15462 10362
rect 15514 10310 15520 10362
rect 552 10288 15520 10310
rect 552 9818 15364 9840
rect 552 9766 2249 9818
rect 2301 9766 2313 9818
rect 2365 9766 2377 9818
rect 2429 9766 2441 9818
rect 2493 9766 2505 9818
rect 2557 9766 5951 9818
rect 6003 9766 6015 9818
rect 6067 9766 6079 9818
rect 6131 9766 6143 9818
rect 6195 9766 6207 9818
rect 6259 9766 9653 9818
rect 9705 9766 9717 9818
rect 9769 9766 9781 9818
rect 9833 9766 9845 9818
rect 9897 9766 9909 9818
rect 9961 9766 13355 9818
rect 13407 9766 13419 9818
rect 13471 9766 13483 9818
rect 13535 9766 13547 9818
rect 13599 9766 13611 9818
rect 13663 9766 15364 9818
rect 552 9744 15364 9766
rect 552 9274 15520 9296
rect 552 9222 4100 9274
rect 4152 9222 4164 9274
rect 4216 9222 4228 9274
rect 4280 9222 4292 9274
rect 4344 9222 4356 9274
rect 4408 9222 7802 9274
rect 7854 9222 7866 9274
rect 7918 9222 7930 9274
rect 7982 9222 7994 9274
rect 8046 9222 8058 9274
rect 8110 9222 11504 9274
rect 11556 9222 11568 9274
rect 11620 9222 11632 9274
rect 11684 9222 11696 9274
rect 11748 9222 11760 9274
rect 11812 9222 15206 9274
rect 15258 9222 15270 9274
rect 15322 9222 15334 9274
rect 15386 9222 15398 9274
rect 15450 9222 15462 9274
rect 15514 9222 15520 9274
rect 552 9200 15520 9222
rect 552 8730 15364 8752
rect 552 8678 2249 8730
rect 2301 8678 2313 8730
rect 2365 8678 2377 8730
rect 2429 8678 2441 8730
rect 2493 8678 2505 8730
rect 2557 8678 5951 8730
rect 6003 8678 6015 8730
rect 6067 8678 6079 8730
rect 6131 8678 6143 8730
rect 6195 8678 6207 8730
rect 6259 8678 9653 8730
rect 9705 8678 9717 8730
rect 9769 8678 9781 8730
rect 9833 8678 9845 8730
rect 9897 8678 9909 8730
rect 9961 8678 13355 8730
rect 13407 8678 13419 8730
rect 13471 8678 13483 8730
rect 13535 8678 13547 8730
rect 13599 8678 13611 8730
rect 13663 8678 15364 8730
rect 552 8656 15364 8678
rect 552 8186 15520 8208
rect 552 8134 4100 8186
rect 4152 8134 4164 8186
rect 4216 8134 4228 8186
rect 4280 8134 4292 8186
rect 4344 8134 4356 8186
rect 4408 8134 7802 8186
rect 7854 8134 7866 8186
rect 7918 8134 7930 8186
rect 7982 8134 7994 8186
rect 8046 8134 8058 8186
rect 8110 8134 11504 8186
rect 11556 8134 11568 8186
rect 11620 8134 11632 8186
rect 11684 8134 11696 8186
rect 11748 8134 11760 8186
rect 11812 8134 15206 8186
rect 15258 8134 15270 8186
rect 15322 8134 15334 8186
rect 15386 8134 15398 8186
rect 15450 8134 15462 8186
rect 15514 8134 15520 8186
rect 552 8112 15520 8134
rect 552 7642 15364 7664
rect 552 7590 2249 7642
rect 2301 7590 2313 7642
rect 2365 7590 2377 7642
rect 2429 7590 2441 7642
rect 2493 7590 2505 7642
rect 2557 7590 5951 7642
rect 6003 7590 6015 7642
rect 6067 7590 6079 7642
rect 6131 7590 6143 7642
rect 6195 7590 6207 7642
rect 6259 7590 9653 7642
rect 9705 7590 9717 7642
rect 9769 7590 9781 7642
rect 9833 7590 9845 7642
rect 9897 7590 9909 7642
rect 9961 7590 13355 7642
rect 13407 7590 13419 7642
rect 13471 7590 13483 7642
rect 13535 7590 13547 7642
rect 13599 7590 13611 7642
rect 13663 7590 15364 7642
rect 552 7568 15364 7590
rect 552 7098 15520 7120
rect 552 7046 4100 7098
rect 4152 7046 4164 7098
rect 4216 7046 4228 7098
rect 4280 7046 4292 7098
rect 4344 7046 4356 7098
rect 4408 7046 7802 7098
rect 7854 7046 7866 7098
rect 7918 7046 7930 7098
rect 7982 7046 7994 7098
rect 8046 7046 8058 7098
rect 8110 7046 11504 7098
rect 11556 7046 11568 7098
rect 11620 7046 11632 7098
rect 11684 7046 11696 7098
rect 11748 7046 11760 7098
rect 11812 7046 15206 7098
rect 15258 7046 15270 7098
rect 15322 7046 15334 7098
rect 15386 7046 15398 7098
rect 15450 7046 15462 7098
rect 15514 7046 15520 7098
rect 552 7024 15520 7046
rect 552 6554 15364 6576
rect 552 6502 2249 6554
rect 2301 6502 2313 6554
rect 2365 6502 2377 6554
rect 2429 6502 2441 6554
rect 2493 6502 2505 6554
rect 2557 6502 5951 6554
rect 6003 6502 6015 6554
rect 6067 6502 6079 6554
rect 6131 6502 6143 6554
rect 6195 6502 6207 6554
rect 6259 6502 9653 6554
rect 9705 6502 9717 6554
rect 9769 6502 9781 6554
rect 9833 6502 9845 6554
rect 9897 6502 9909 6554
rect 9961 6502 13355 6554
rect 13407 6502 13419 6554
rect 13471 6502 13483 6554
rect 13535 6502 13547 6554
rect 13599 6502 13611 6554
rect 13663 6502 15364 6554
rect 552 6480 15364 6502
rect 552 6010 15520 6032
rect 552 5958 4100 6010
rect 4152 5958 4164 6010
rect 4216 5958 4228 6010
rect 4280 5958 4292 6010
rect 4344 5958 4356 6010
rect 4408 5958 7802 6010
rect 7854 5958 7866 6010
rect 7918 5958 7930 6010
rect 7982 5958 7994 6010
rect 8046 5958 8058 6010
rect 8110 5958 11504 6010
rect 11556 5958 11568 6010
rect 11620 5958 11632 6010
rect 11684 5958 11696 6010
rect 11748 5958 11760 6010
rect 11812 5958 15206 6010
rect 15258 5958 15270 6010
rect 15322 5958 15334 6010
rect 15386 5958 15398 6010
rect 15450 5958 15462 6010
rect 15514 5958 15520 6010
rect 552 5936 15520 5958
rect 552 5466 15364 5488
rect 552 5414 2249 5466
rect 2301 5414 2313 5466
rect 2365 5414 2377 5466
rect 2429 5414 2441 5466
rect 2493 5414 2505 5466
rect 2557 5414 5951 5466
rect 6003 5414 6015 5466
rect 6067 5414 6079 5466
rect 6131 5414 6143 5466
rect 6195 5414 6207 5466
rect 6259 5414 9653 5466
rect 9705 5414 9717 5466
rect 9769 5414 9781 5466
rect 9833 5414 9845 5466
rect 9897 5414 9909 5466
rect 9961 5414 13355 5466
rect 13407 5414 13419 5466
rect 13471 5414 13483 5466
rect 13535 5414 13547 5466
rect 13599 5414 13611 5466
rect 13663 5414 15364 5466
rect 552 5392 15364 5414
rect 552 4922 15520 4944
rect 552 4870 4100 4922
rect 4152 4870 4164 4922
rect 4216 4870 4228 4922
rect 4280 4870 4292 4922
rect 4344 4870 4356 4922
rect 4408 4870 7802 4922
rect 7854 4870 7866 4922
rect 7918 4870 7930 4922
rect 7982 4870 7994 4922
rect 8046 4870 8058 4922
rect 8110 4870 11504 4922
rect 11556 4870 11568 4922
rect 11620 4870 11632 4922
rect 11684 4870 11696 4922
rect 11748 4870 11760 4922
rect 11812 4870 15206 4922
rect 15258 4870 15270 4922
rect 15322 4870 15334 4922
rect 15386 4870 15398 4922
rect 15450 4870 15462 4922
rect 15514 4870 15520 4922
rect 552 4848 15520 4870
rect 11330 4700 11336 4752
rect 11388 4700 11394 4752
rect 11238 4428 11244 4480
rect 11296 4428 11302 4480
rect 552 4378 15364 4400
rect 552 4326 2249 4378
rect 2301 4326 2313 4378
rect 2365 4326 2377 4378
rect 2429 4326 2441 4378
rect 2493 4326 2505 4378
rect 2557 4326 5951 4378
rect 6003 4326 6015 4378
rect 6067 4326 6079 4378
rect 6131 4326 6143 4378
rect 6195 4326 6207 4378
rect 6259 4326 9653 4378
rect 9705 4326 9717 4378
rect 9769 4326 9781 4378
rect 9833 4326 9845 4378
rect 9897 4326 9909 4378
rect 9961 4326 13355 4378
rect 13407 4326 13419 4378
rect 13471 4326 13483 4378
rect 13535 4326 13547 4378
rect 13599 4326 13611 4378
rect 13663 4326 15364 4378
rect 552 4304 15364 4326
rect 552 3834 15520 3856
rect 552 3782 4100 3834
rect 4152 3782 4164 3834
rect 4216 3782 4228 3834
rect 4280 3782 4292 3834
rect 4344 3782 4356 3834
rect 4408 3782 7802 3834
rect 7854 3782 7866 3834
rect 7918 3782 7930 3834
rect 7982 3782 7994 3834
rect 8046 3782 8058 3834
rect 8110 3782 11504 3834
rect 11556 3782 11568 3834
rect 11620 3782 11632 3834
rect 11684 3782 11696 3834
rect 11748 3782 11760 3834
rect 11812 3782 15206 3834
rect 15258 3782 15270 3834
rect 15322 3782 15334 3834
rect 15386 3782 15398 3834
rect 15450 3782 15462 3834
rect 15514 3782 15520 3834
rect 552 3760 15520 3782
rect 552 3290 15364 3312
rect 552 3238 2249 3290
rect 2301 3238 2313 3290
rect 2365 3238 2377 3290
rect 2429 3238 2441 3290
rect 2493 3238 2505 3290
rect 2557 3238 5951 3290
rect 6003 3238 6015 3290
rect 6067 3238 6079 3290
rect 6131 3238 6143 3290
rect 6195 3238 6207 3290
rect 6259 3238 9653 3290
rect 9705 3238 9717 3290
rect 9769 3238 9781 3290
rect 9833 3238 9845 3290
rect 9897 3238 9909 3290
rect 9961 3238 13355 3290
rect 13407 3238 13419 3290
rect 13471 3238 13483 3290
rect 13535 3238 13547 3290
rect 13599 3238 13611 3290
rect 13663 3238 15364 3290
rect 552 3216 15364 3238
rect 552 2746 15520 2768
rect 552 2694 4100 2746
rect 4152 2694 4164 2746
rect 4216 2694 4228 2746
rect 4280 2694 4292 2746
rect 4344 2694 4356 2746
rect 4408 2694 7802 2746
rect 7854 2694 7866 2746
rect 7918 2694 7930 2746
rect 7982 2694 7994 2746
rect 8046 2694 8058 2746
rect 8110 2694 11504 2746
rect 11556 2694 11568 2746
rect 11620 2694 11632 2746
rect 11684 2694 11696 2746
rect 11748 2694 11760 2746
rect 11812 2694 15206 2746
rect 15258 2694 15270 2746
rect 15322 2694 15334 2746
rect 15386 2694 15398 2746
rect 15450 2694 15462 2746
rect 15514 2694 15520 2746
rect 552 2672 15520 2694
rect 552 2202 15364 2224
rect 552 2150 2249 2202
rect 2301 2150 2313 2202
rect 2365 2150 2377 2202
rect 2429 2150 2441 2202
rect 2493 2150 2505 2202
rect 2557 2150 5951 2202
rect 6003 2150 6015 2202
rect 6067 2150 6079 2202
rect 6131 2150 6143 2202
rect 6195 2150 6207 2202
rect 6259 2150 9653 2202
rect 9705 2150 9717 2202
rect 9769 2150 9781 2202
rect 9833 2150 9845 2202
rect 9897 2150 9909 2202
rect 9961 2150 13355 2202
rect 13407 2150 13419 2202
rect 13471 2150 13483 2202
rect 13535 2150 13547 2202
rect 13599 2150 13611 2202
rect 13663 2150 15364 2202
rect 552 2128 15364 2150
rect 552 1658 15520 1680
rect 552 1606 4100 1658
rect 4152 1606 4164 1658
rect 4216 1606 4228 1658
rect 4280 1606 4292 1658
rect 4344 1606 4356 1658
rect 4408 1606 7802 1658
rect 7854 1606 7866 1658
rect 7918 1606 7930 1658
rect 7982 1606 7994 1658
rect 8046 1606 8058 1658
rect 8110 1606 11504 1658
rect 11556 1606 11568 1658
rect 11620 1606 11632 1658
rect 11684 1606 11696 1658
rect 11748 1606 11760 1658
rect 11812 1606 15206 1658
rect 15258 1606 15270 1658
rect 15322 1606 15334 1658
rect 15386 1606 15398 1658
rect 15450 1606 15462 1658
rect 15514 1606 15520 1658
rect 552 1584 15520 1606
rect 552 1114 15364 1136
rect 552 1062 2249 1114
rect 2301 1062 2313 1114
rect 2365 1062 2377 1114
rect 2429 1062 2441 1114
rect 2493 1062 2505 1114
rect 2557 1062 5951 1114
rect 6003 1062 6015 1114
rect 6067 1062 6079 1114
rect 6131 1062 6143 1114
rect 6195 1062 6207 1114
rect 6259 1062 9653 1114
rect 9705 1062 9717 1114
rect 9769 1062 9781 1114
rect 9833 1062 9845 1114
rect 9897 1062 9909 1114
rect 9961 1062 13355 1114
rect 13407 1062 13419 1114
rect 13471 1062 13483 1114
rect 13535 1062 13547 1114
rect 13599 1062 13611 1114
rect 13663 1062 15364 1114
rect 552 1040 15364 1062
rect 552 570 15520 592
rect 552 518 4100 570
rect 4152 518 4164 570
rect 4216 518 4228 570
rect 4280 518 4292 570
rect 4344 518 4356 570
rect 4408 518 7802 570
rect 7854 518 7866 570
rect 7918 518 7930 570
rect 7982 518 7994 570
rect 8046 518 8058 570
rect 8110 518 11504 570
rect 11556 518 11568 570
rect 11620 518 11632 570
rect 11684 518 11696 570
rect 11748 518 11760 570
rect 11812 518 15206 570
rect 15258 518 15270 570
rect 15322 518 15334 570
rect 15386 518 15398 570
rect 15450 518 15462 570
rect 15514 518 15520 570
rect 552 496 15520 518
<< via1 >>
rect 2249 15206 2301 15258
rect 2313 15206 2365 15258
rect 2377 15206 2429 15258
rect 2441 15206 2493 15258
rect 2505 15206 2557 15258
rect 5951 15206 6003 15258
rect 6015 15206 6067 15258
rect 6079 15206 6131 15258
rect 6143 15206 6195 15258
rect 6207 15206 6259 15258
rect 9653 15206 9705 15258
rect 9717 15206 9769 15258
rect 9781 15206 9833 15258
rect 9845 15206 9897 15258
rect 9909 15206 9961 15258
rect 13355 15206 13407 15258
rect 13419 15206 13471 15258
rect 13483 15206 13535 15258
rect 13547 15206 13599 15258
rect 13611 15206 13663 15258
rect 9404 15147 9456 15156
rect 9404 15113 9413 15147
rect 9413 15113 9447 15147
rect 9447 15113 9456 15147
rect 9404 15104 9456 15113
rect 1216 14900 1268 14952
rect 3148 14900 3200 14952
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 3976 14764 4028 14816
rect 4528 14832 4580 14884
rect 10968 15011 11020 15020
rect 10968 14977 10977 15011
rect 10977 14977 11011 15011
rect 11011 14977 11020 15011
rect 10968 14968 11020 14977
rect 5080 14900 5132 14952
rect 6552 14900 6604 14952
rect 7104 14900 7156 14952
rect 8760 14900 8812 14952
rect 5632 14832 5684 14884
rect 9680 14943 9732 14952
rect 9680 14909 9689 14943
rect 9689 14909 9723 14943
rect 9723 14909 9732 14943
rect 9680 14900 9732 14909
rect 12440 14900 12492 14952
rect 12808 14900 12860 14952
rect 11980 14832 12032 14884
rect 4436 14807 4488 14816
rect 4436 14773 4445 14807
rect 4445 14773 4479 14807
rect 4479 14773 4488 14807
rect 4436 14764 4488 14773
rect 4712 14764 4764 14816
rect 6276 14807 6328 14816
rect 6276 14773 6285 14807
rect 6285 14773 6319 14807
rect 6319 14773 6328 14807
rect 6276 14764 6328 14773
rect 8760 14807 8812 14816
rect 8760 14773 8769 14807
rect 8769 14773 8803 14807
rect 8803 14773 8812 14807
rect 8760 14764 8812 14773
rect 9312 14764 9364 14816
rect 10324 14807 10376 14816
rect 10324 14773 10333 14807
rect 10333 14773 10367 14807
rect 10367 14773 10376 14807
rect 10324 14764 10376 14773
rect 10416 14764 10468 14816
rect 11888 14807 11940 14816
rect 11888 14773 11897 14807
rect 11897 14773 11931 14807
rect 11931 14773 11940 14807
rect 11888 14764 11940 14773
rect 13084 14807 13136 14816
rect 13084 14773 13093 14807
rect 13093 14773 13127 14807
rect 13127 14773 13136 14807
rect 13084 14764 13136 14773
rect 4100 14662 4152 14714
rect 4164 14662 4216 14714
rect 4228 14662 4280 14714
rect 4292 14662 4344 14714
rect 4356 14662 4408 14714
rect 7802 14662 7854 14714
rect 7866 14662 7918 14714
rect 7930 14662 7982 14714
rect 7994 14662 8046 14714
rect 8058 14662 8110 14714
rect 11504 14662 11556 14714
rect 11568 14662 11620 14714
rect 11632 14662 11684 14714
rect 11696 14662 11748 14714
rect 11760 14662 11812 14714
rect 15206 14662 15258 14714
rect 15270 14662 15322 14714
rect 15334 14662 15386 14714
rect 15398 14662 15450 14714
rect 15462 14662 15514 14714
rect 1492 14560 1544 14612
rect 3976 14560 4028 14612
rect 8668 14560 8720 14612
rect 8760 14560 8812 14612
rect 4528 14492 4580 14544
rect 4436 14467 4488 14476
rect 4436 14433 4445 14467
rect 4445 14433 4479 14467
rect 4479 14433 4488 14467
rect 4436 14424 4488 14433
rect 4620 14467 4672 14476
rect 4620 14433 4629 14467
rect 4629 14433 4663 14467
rect 4663 14433 4672 14467
rect 4620 14424 4672 14433
rect 4528 14331 4580 14340
rect 4528 14297 4537 14331
rect 4537 14297 4571 14331
rect 4571 14297 4580 14331
rect 4528 14288 4580 14297
rect 5356 14467 5408 14476
rect 5356 14433 5365 14467
rect 5365 14433 5399 14467
rect 5399 14433 5408 14467
rect 5356 14424 5408 14433
rect 5448 14467 5500 14476
rect 5448 14433 5457 14467
rect 5457 14433 5491 14467
rect 5491 14433 5500 14467
rect 5448 14424 5500 14433
rect 5172 14288 5224 14340
rect 5632 14331 5684 14340
rect 5632 14297 5641 14331
rect 5641 14297 5675 14331
rect 5675 14297 5684 14331
rect 5632 14288 5684 14297
rect 7104 14424 7156 14476
rect 7564 14424 7616 14476
rect 9404 14492 9456 14544
rect 8392 14424 8444 14476
rect 6368 14356 6420 14408
rect 6552 14288 6604 14340
rect 9680 14560 9732 14612
rect 10324 14560 10376 14612
rect 13820 14560 13872 14612
rect 13084 14424 13136 14476
rect 11336 14356 11388 14408
rect 11796 14356 11848 14408
rect 5816 14220 5868 14272
rect 7380 14220 7432 14272
rect 9312 14220 9364 14272
rect 9496 14220 9548 14272
rect 10416 14220 10468 14272
rect 13268 14263 13320 14272
rect 13268 14229 13277 14263
rect 13277 14229 13311 14263
rect 13311 14229 13320 14263
rect 13268 14220 13320 14229
rect 2249 14118 2301 14170
rect 2313 14118 2365 14170
rect 2377 14118 2429 14170
rect 2441 14118 2493 14170
rect 2505 14118 2557 14170
rect 5951 14118 6003 14170
rect 6015 14118 6067 14170
rect 6079 14118 6131 14170
rect 6143 14118 6195 14170
rect 6207 14118 6259 14170
rect 9653 14118 9705 14170
rect 9717 14118 9769 14170
rect 9781 14118 9833 14170
rect 9845 14118 9897 14170
rect 9909 14118 9961 14170
rect 13355 14118 13407 14170
rect 13419 14118 13471 14170
rect 13483 14118 13535 14170
rect 13547 14118 13599 14170
rect 13611 14118 13663 14170
rect 3976 14016 4028 14068
rect 4528 14016 4580 14068
rect 5448 14016 5500 14068
rect 6276 14016 6328 14068
rect 5172 13880 5224 13932
rect 4712 13812 4764 13864
rect 5264 13812 5316 13864
rect 5356 13676 5408 13728
rect 5816 13719 5868 13728
rect 5816 13685 5825 13719
rect 5825 13685 5859 13719
rect 5859 13685 5868 13719
rect 5816 13676 5868 13685
rect 6368 13812 6420 13864
rect 7196 14016 7248 14068
rect 7380 13948 7432 14000
rect 7564 14016 7616 14068
rect 8392 14059 8444 14068
rect 8392 14025 8401 14059
rect 8401 14025 8435 14059
rect 8435 14025 8444 14059
rect 8392 14016 8444 14025
rect 9404 14016 9456 14068
rect 10416 14016 10468 14068
rect 11428 14016 11480 14068
rect 12440 14016 12492 14068
rect 6736 13676 6788 13728
rect 8208 13812 8260 13864
rect 8668 13812 8720 13864
rect 9496 13880 9548 13932
rect 14740 13948 14792 14000
rect 11980 13880 12032 13932
rect 12440 13923 12492 13932
rect 12440 13889 12449 13923
rect 12449 13889 12483 13923
rect 12483 13889 12492 13923
rect 12440 13880 12492 13889
rect 11888 13812 11940 13864
rect 13268 13880 13320 13932
rect 9772 13744 9824 13796
rect 11244 13744 11296 13796
rect 10048 13676 10100 13728
rect 12256 13719 12308 13728
rect 12256 13685 12265 13719
rect 12265 13685 12299 13719
rect 12299 13685 12308 13719
rect 12256 13676 12308 13685
rect 13268 13676 13320 13728
rect 4100 13574 4152 13626
rect 4164 13574 4216 13626
rect 4228 13574 4280 13626
rect 4292 13574 4344 13626
rect 4356 13574 4408 13626
rect 7802 13574 7854 13626
rect 7866 13574 7918 13626
rect 7930 13574 7982 13626
rect 7994 13574 8046 13626
rect 8058 13574 8110 13626
rect 11504 13574 11556 13626
rect 11568 13574 11620 13626
rect 11632 13574 11684 13626
rect 11696 13574 11748 13626
rect 11760 13574 11812 13626
rect 15206 13574 15258 13626
rect 15270 13574 15322 13626
rect 15334 13574 15386 13626
rect 15398 13574 15450 13626
rect 15462 13574 15514 13626
rect 4620 13472 4672 13524
rect 11244 13472 11296 13524
rect 12256 13472 12308 13524
rect 10048 13404 10100 13456
rect 5356 13336 5408 13388
rect 7380 13336 7432 13388
rect 9772 13336 9824 13388
rect 10876 13336 10928 13388
rect 5172 13311 5224 13320
rect 5172 13277 5181 13311
rect 5181 13277 5215 13311
rect 5215 13277 5224 13311
rect 5172 13268 5224 13277
rect 4804 13200 4856 13252
rect 11888 13268 11940 13320
rect 10876 13200 10928 13252
rect 7104 13132 7156 13184
rect 7840 13175 7892 13184
rect 7840 13141 7849 13175
rect 7849 13141 7883 13175
rect 7883 13141 7892 13175
rect 7840 13132 7892 13141
rect 12256 13175 12308 13184
rect 12256 13141 12265 13175
rect 12265 13141 12299 13175
rect 12299 13141 12308 13175
rect 12256 13132 12308 13141
rect 2249 13030 2301 13082
rect 2313 13030 2365 13082
rect 2377 13030 2429 13082
rect 2441 13030 2493 13082
rect 2505 13030 2557 13082
rect 5951 13030 6003 13082
rect 6015 13030 6067 13082
rect 6079 13030 6131 13082
rect 6143 13030 6195 13082
rect 6207 13030 6259 13082
rect 9653 13030 9705 13082
rect 9717 13030 9769 13082
rect 9781 13030 9833 13082
rect 9845 13030 9897 13082
rect 9909 13030 9961 13082
rect 13355 13030 13407 13082
rect 13419 13030 13471 13082
rect 13483 13030 13535 13082
rect 13547 13030 13599 13082
rect 13611 13030 13663 13082
rect 4712 12928 4764 12980
rect 4804 12971 4856 12980
rect 4804 12937 4813 12971
rect 4813 12937 4847 12971
rect 4847 12937 4856 12971
rect 4804 12928 4856 12937
rect 5172 12928 5224 12980
rect 6736 12971 6788 12980
rect 6736 12937 6745 12971
rect 6745 12937 6779 12971
rect 6779 12937 6788 12971
rect 6736 12928 6788 12937
rect 10876 12928 10928 12980
rect 7104 12792 7156 12844
rect 5264 12724 5316 12776
rect 5908 12767 5960 12776
rect 5908 12733 5917 12767
rect 5917 12733 5951 12767
rect 5951 12733 5960 12767
rect 5908 12724 5960 12733
rect 7012 12724 7064 12776
rect 11336 12724 11388 12776
rect 12256 12724 12308 12776
rect 6736 12588 6788 12640
rect 7840 12699 7892 12708
rect 7840 12665 7858 12699
rect 7858 12665 7892 12699
rect 7840 12656 7892 12665
rect 9404 12656 9456 12708
rect 13268 12656 13320 12708
rect 8392 12631 8444 12640
rect 8392 12597 8401 12631
rect 8401 12597 8435 12631
rect 8435 12597 8444 12631
rect 8392 12588 8444 12597
rect 4100 12486 4152 12538
rect 4164 12486 4216 12538
rect 4228 12486 4280 12538
rect 4292 12486 4344 12538
rect 4356 12486 4408 12538
rect 7802 12486 7854 12538
rect 7866 12486 7918 12538
rect 7930 12486 7982 12538
rect 7994 12486 8046 12538
rect 8058 12486 8110 12538
rect 11504 12486 11556 12538
rect 11568 12486 11620 12538
rect 11632 12486 11684 12538
rect 11696 12486 11748 12538
rect 11760 12486 11812 12538
rect 15206 12486 15258 12538
rect 15270 12486 15322 12538
rect 15334 12486 15386 12538
rect 15398 12486 15450 12538
rect 15462 12486 15514 12538
rect 4712 12384 4764 12436
rect 5356 12427 5408 12436
rect 5356 12393 5365 12427
rect 5365 12393 5399 12427
rect 5399 12393 5408 12427
rect 5356 12384 5408 12393
rect 7104 12384 7156 12436
rect 7196 12427 7248 12436
rect 7196 12393 7205 12427
rect 7205 12393 7239 12427
rect 7239 12393 7248 12427
rect 7196 12384 7248 12393
rect 8208 12384 8260 12436
rect 8392 12248 8444 12300
rect 9404 12384 9456 12436
rect 9312 12248 9364 12300
rect 13820 12248 13872 12300
rect 5816 12044 5868 12096
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 14740 12087 14792 12096
rect 14740 12053 14749 12087
rect 14749 12053 14783 12087
rect 14783 12053 14792 12087
rect 14740 12044 14792 12053
rect 2249 11942 2301 11994
rect 2313 11942 2365 11994
rect 2377 11942 2429 11994
rect 2441 11942 2493 11994
rect 2505 11942 2557 11994
rect 5951 11942 6003 11994
rect 6015 11942 6067 11994
rect 6079 11942 6131 11994
rect 6143 11942 6195 11994
rect 6207 11942 6259 11994
rect 9653 11942 9705 11994
rect 9717 11942 9769 11994
rect 9781 11942 9833 11994
rect 9845 11942 9897 11994
rect 9909 11942 9961 11994
rect 13355 11942 13407 11994
rect 13419 11942 13471 11994
rect 13483 11942 13535 11994
rect 13547 11942 13599 11994
rect 13611 11942 13663 11994
rect 4100 11398 4152 11450
rect 4164 11398 4216 11450
rect 4228 11398 4280 11450
rect 4292 11398 4344 11450
rect 4356 11398 4408 11450
rect 7802 11398 7854 11450
rect 7866 11398 7918 11450
rect 7930 11398 7982 11450
rect 7994 11398 8046 11450
rect 8058 11398 8110 11450
rect 11504 11398 11556 11450
rect 11568 11398 11620 11450
rect 11632 11398 11684 11450
rect 11696 11398 11748 11450
rect 11760 11398 11812 11450
rect 15206 11398 15258 11450
rect 15270 11398 15322 11450
rect 15334 11398 15386 11450
rect 15398 11398 15450 11450
rect 15462 11398 15514 11450
rect 2249 10854 2301 10906
rect 2313 10854 2365 10906
rect 2377 10854 2429 10906
rect 2441 10854 2493 10906
rect 2505 10854 2557 10906
rect 5951 10854 6003 10906
rect 6015 10854 6067 10906
rect 6079 10854 6131 10906
rect 6143 10854 6195 10906
rect 6207 10854 6259 10906
rect 9653 10854 9705 10906
rect 9717 10854 9769 10906
rect 9781 10854 9833 10906
rect 9845 10854 9897 10906
rect 9909 10854 9961 10906
rect 13355 10854 13407 10906
rect 13419 10854 13471 10906
rect 13483 10854 13535 10906
rect 13547 10854 13599 10906
rect 13611 10854 13663 10906
rect 4100 10310 4152 10362
rect 4164 10310 4216 10362
rect 4228 10310 4280 10362
rect 4292 10310 4344 10362
rect 4356 10310 4408 10362
rect 7802 10310 7854 10362
rect 7866 10310 7918 10362
rect 7930 10310 7982 10362
rect 7994 10310 8046 10362
rect 8058 10310 8110 10362
rect 11504 10310 11556 10362
rect 11568 10310 11620 10362
rect 11632 10310 11684 10362
rect 11696 10310 11748 10362
rect 11760 10310 11812 10362
rect 15206 10310 15258 10362
rect 15270 10310 15322 10362
rect 15334 10310 15386 10362
rect 15398 10310 15450 10362
rect 15462 10310 15514 10362
rect 2249 9766 2301 9818
rect 2313 9766 2365 9818
rect 2377 9766 2429 9818
rect 2441 9766 2493 9818
rect 2505 9766 2557 9818
rect 5951 9766 6003 9818
rect 6015 9766 6067 9818
rect 6079 9766 6131 9818
rect 6143 9766 6195 9818
rect 6207 9766 6259 9818
rect 9653 9766 9705 9818
rect 9717 9766 9769 9818
rect 9781 9766 9833 9818
rect 9845 9766 9897 9818
rect 9909 9766 9961 9818
rect 13355 9766 13407 9818
rect 13419 9766 13471 9818
rect 13483 9766 13535 9818
rect 13547 9766 13599 9818
rect 13611 9766 13663 9818
rect 4100 9222 4152 9274
rect 4164 9222 4216 9274
rect 4228 9222 4280 9274
rect 4292 9222 4344 9274
rect 4356 9222 4408 9274
rect 7802 9222 7854 9274
rect 7866 9222 7918 9274
rect 7930 9222 7982 9274
rect 7994 9222 8046 9274
rect 8058 9222 8110 9274
rect 11504 9222 11556 9274
rect 11568 9222 11620 9274
rect 11632 9222 11684 9274
rect 11696 9222 11748 9274
rect 11760 9222 11812 9274
rect 15206 9222 15258 9274
rect 15270 9222 15322 9274
rect 15334 9222 15386 9274
rect 15398 9222 15450 9274
rect 15462 9222 15514 9274
rect 2249 8678 2301 8730
rect 2313 8678 2365 8730
rect 2377 8678 2429 8730
rect 2441 8678 2493 8730
rect 2505 8678 2557 8730
rect 5951 8678 6003 8730
rect 6015 8678 6067 8730
rect 6079 8678 6131 8730
rect 6143 8678 6195 8730
rect 6207 8678 6259 8730
rect 9653 8678 9705 8730
rect 9717 8678 9769 8730
rect 9781 8678 9833 8730
rect 9845 8678 9897 8730
rect 9909 8678 9961 8730
rect 13355 8678 13407 8730
rect 13419 8678 13471 8730
rect 13483 8678 13535 8730
rect 13547 8678 13599 8730
rect 13611 8678 13663 8730
rect 4100 8134 4152 8186
rect 4164 8134 4216 8186
rect 4228 8134 4280 8186
rect 4292 8134 4344 8186
rect 4356 8134 4408 8186
rect 7802 8134 7854 8186
rect 7866 8134 7918 8186
rect 7930 8134 7982 8186
rect 7994 8134 8046 8186
rect 8058 8134 8110 8186
rect 11504 8134 11556 8186
rect 11568 8134 11620 8186
rect 11632 8134 11684 8186
rect 11696 8134 11748 8186
rect 11760 8134 11812 8186
rect 15206 8134 15258 8186
rect 15270 8134 15322 8186
rect 15334 8134 15386 8186
rect 15398 8134 15450 8186
rect 15462 8134 15514 8186
rect 2249 7590 2301 7642
rect 2313 7590 2365 7642
rect 2377 7590 2429 7642
rect 2441 7590 2493 7642
rect 2505 7590 2557 7642
rect 5951 7590 6003 7642
rect 6015 7590 6067 7642
rect 6079 7590 6131 7642
rect 6143 7590 6195 7642
rect 6207 7590 6259 7642
rect 9653 7590 9705 7642
rect 9717 7590 9769 7642
rect 9781 7590 9833 7642
rect 9845 7590 9897 7642
rect 9909 7590 9961 7642
rect 13355 7590 13407 7642
rect 13419 7590 13471 7642
rect 13483 7590 13535 7642
rect 13547 7590 13599 7642
rect 13611 7590 13663 7642
rect 4100 7046 4152 7098
rect 4164 7046 4216 7098
rect 4228 7046 4280 7098
rect 4292 7046 4344 7098
rect 4356 7046 4408 7098
rect 7802 7046 7854 7098
rect 7866 7046 7918 7098
rect 7930 7046 7982 7098
rect 7994 7046 8046 7098
rect 8058 7046 8110 7098
rect 11504 7046 11556 7098
rect 11568 7046 11620 7098
rect 11632 7046 11684 7098
rect 11696 7046 11748 7098
rect 11760 7046 11812 7098
rect 15206 7046 15258 7098
rect 15270 7046 15322 7098
rect 15334 7046 15386 7098
rect 15398 7046 15450 7098
rect 15462 7046 15514 7098
rect 2249 6502 2301 6554
rect 2313 6502 2365 6554
rect 2377 6502 2429 6554
rect 2441 6502 2493 6554
rect 2505 6502 2557 6554
rect 5951 6502 6003 6554
rect 6015 6502 6067 6554
rect 6079 6502 6131 6554
rect 6143 6502 6195 6554
rect 6207 6502 6259 6554
rect 9653 6502 9705 6554
rect 9717 6502 9769 6554
rect 9781 6502 9833 6554
rect 9845 6502 9897 6554
rect 9909 6502 9961 6554
rect 13355 6502 13407 6554
rect 13419 6502 13471 6554
rect 13483 6502 13535 6554
rect 13547 6502 13599 6554
rect 13611 6502 13663 6554
rect 4100 5958 4152 6010
rect 4164 5958 4216 6010
rect 4228 5958 4280 6010
rect 4292 5958 4344 6010
rect 4356 5958 4408 6010
rect 7802 5958 7854 6010
rect 7866 5958 7918 6010
rect 7930 5958 7982 6010
rect 7994 5958 8046 6010
rect 8058 5958 8110 6010
rect 11504 5958 11556 6010
rect 11568 5958 11620 6010
rect 11632 5958 11684 6010
rect 11696 5958 11748 6010
rect 11760 5958 11812 6010
rect 15206 5958 15258 6010
rect 15270 5958 15322 6010
rect 15334 5958 15386 6010
rect 15398 5958 15450 6010
rect 15462 5958 15514 6010
rect 2249 5414 2301 5466
rect 2313 5414 2365 5466
rect 2377 5414 2429 5466
rect 2441 5414 2493 5466
rect 2505 5414 2557 5466
rect 5951 5414 6003 5466
rect 6015 5414 6067 5466
rect 6079 5414 6131 5466
rect 6143 5414 6195 5466
rect 6207 5414 6259 5466
rect 9653 5414 9705 5466
rect 9717 5414 9769 5466
rect 9781 5414 9833 5466
rect 9845 5414 9897 5466
rect 9909 5414 9961 5466
rect 13355 5414 13407 5466
rect 13419 5414 13471 5466
rect 13483 5414 13535 5466
rect 13547 5414 13599 5466
rect 13611 5414 13663 5466
rect 4100 4870 4152 4922
rect 4164 4870 4216 4922
rect 4228 4870 4280 4922
rect 4292 4870 4344 4922
rect 4356 4870 4408 4922
rect 7802 4870 7854 4922
rect 7866 4870 7918 4922
rect 7930 4870 7982 4922
rect 7994 4870 8046 4922
rect 8058 4870 8110 4922
rect 11504 4870 11556 4922
rect 11568 4870 11620 4922
rect 11632 4870 11684 4922
rect 11696 4870 11748 4922
rect 11760 4870 11812 4922
rect 15206 4870 15258 4922
rect 15270 4870 15322 4922
rect 15334 4870 15386 4922
rect 15398 4870 15450 4922
rect 15462 4870 15514 4922
rect 11336 4743 11388 4752
rect 11336 4709 11345 4743
rect 11345 4709 11379 4743
rect 11379 4709 11388 4743
rect 11336 4700 11388 4709
rect 11244 4471 11296 4480
rect 11244 4437 11253 4471
rect 11253 4437 11287 4471
rect 11287 4437 11296 4471
rect 11244 4428 11296 4437
rect 2249 4326 2301 4378
rect 2313 4326 2365 4378
rect 2377 4326 2429 4378
rect 2441 4326 2493 4378
rect 2505 4326 2557 4378
rect 5951 4326 6003 4378
rect 6015 4326 6067 4378
rect 6079 4326 6131 4378
rect 6143 4326 6195 4378
rect 6207 4326 6259 4378
rect 9653 4326 9705 4378
rect 9717 4326 9769 4378
rect 9781 4326 9833 4378
rect 9845 4326 9897 4378
rect 9909 4326 9961 4378
rect 13355 4326 13407 4378
rect 13419 4326 13471 4378
rect 13483 4326 13535 4378
rect 13547 4326 13599 4378
rect 13611 4326 13663 4378
rect 4100 3782 4152 3834
rect 4164 3782 4216 3834
rect 4228 3782 4280 3834
rect 4292 3782 4344 3834
rect 4356 3782 4408 3834
rect 7802 3782 7854 3834
rect 7866 3782 7918 3834
rect 7930 3782 7982 3834
rect 7994 3782 8046 3834
rect 8058 3782 8110 3834
rect 11504 3782 11556 3834
rect 11568 3782 11620 3834
rect 11632 3782 11684 3834
rect 11696 3782 11748 3834
rect 11760 3782 11812 3834
rect 15206 3782 15258 3834
rect 15270 3782 15322 3834
rect 15334 3782 15386 3834
rect 15398 3782 15450 3834
rect 15462 3782 15514 3834
rect 2249 3238 2301 3290
rect 2313 3238 2365 3290
rect 2377 3238 2429 3290
rect 2441 3238 2493 3290
rect 2505 3238 2557 3290
rect 5951 3238 6003 3290
rect 6015 3238 6067 3290
rect 6079 3238 6131 3290
rect 6143 3238 6195 3290
rect 6207 3238 6259 3290
rect 9653 3238 9705 3290
rect 9717 3238 9769 3290
rect 9781 3238 9833 3290
rect 9845 3238 9897 3290
rect 9909 3238 9961 3290
rect 13355 3238 13407 3290
rect 13419 3238 13471 3290
rect 13483 3238 13535 3290
rect 13547 3238 13599 3290
rect 13611 3238 13663 3290
rect 4100 2694 4152 2746
rect 4164 2694 4216 2746
rect 4228 2694 4280 2746
rect 4292 2694 4344 2746
rect 4356 2694 4408 2746
rect 7802 2694 7854 2746
rect 7866 2694 7918 2746
rect 7930 2694 7982 2746
rect 7994 2694 8046 2746
rect 8058 2694 8110 2746
rect 11504 2694 11556 2746
rect 11568 2694 11620 2746
rect 11632 2694 11684 2746
rect 11696 2694 11748 2746
rect 11760 2694 11812 2746
rect 15206 2694 15258 2746
rect 15270 2694 15322 2746
rect 15334 2694 15386 2746
rect 15398 2694 15450 2746
rect 15462 2694 15514 2746
rect 2249 2150 2301 2202
rect 2313 2150 2365 2202
rect 2377 2150 2429 2202
rect 2441 2150 2493 2202
rect 2505 2150 2557 2202
rect 5951 2150 6003 2202
rect 6015 2150 6067 2202
rect 6079 2150 6131 2202
rect 6143 2150 6195 2202
rect 6207 2150 6259 2202
rect 9653 2150 9705 2202
rect 9717 2150 9769 2202
rect 9781 2150 9833 2202
rect 9845 2150 9897 2202
rect 9909 2150 9961 2202
rect 13355 2150 13407 2202
rect 13419 2150 13471 2202
rect 13483 2150 13535 2202
rect 13547 2150 13599 2202
rect 13611 2150 13663 2202
rect 4100 1606 4152 1658
rect 4164 1606 4216 1658
rect 4228 1606 4280 1658
rect 4292 1606 4344 1658
rect 4356 1606 4408 1658
rect 7802 1606 7854 1658
rect 7866 1606 7918 1658
rect 7930 1606 7982 1658
rect 7994 1606 8046 1658
rect 8058 1606 8110 1658
rect 11504 1606 11556 1658
rect 11568 1606 11620 1658
rect 11632 1606 11684 1658
rect 11696 1606 11748 1658
rect 11760 1606 11812 1658
rect 15206 1606 15258 1658
rect 15270 1606 15322 1658
rect 15334 1606 15386 1658
rect 15398 1606 15450 1658
rect 15462 1606 15514 1658
rect 2249 1062 2301 1114
rect 2313 1062 2365 1114
rect 2377 1062 2429 1114
rect 2441 1062 2493 1114
rect 2505 1062 2557 1114
rect 5951 1062 6003 1114
rect 6015 1062 6067 1114
rect 6079 1062 6131 1114
rect 6143 1062 6195 1114
rect 6207 1062 6259 1114
rect 9653 1062 9705 1114
rect 9717 1062 9769 1114
rect 9781 1062 9833 1114
rect 9845 1062 9897 1114
rect 9909 1062 9961 1114
rect 13355 1062 13407 1114
rect 13419 1062 13471 1114
rect 13483 1062 13535 1114
rect 13547 1062 13599 1114
rect 13611 1062 13663 1114
rect 4100 518 4152 570
rect 4164 518 4216 570
rect 4228 518 4280 570
rect 4292 518 4344 570
rect 4356 518 4408 570
rect 7802 518 7854 570
rect 7866 518 7918 570
rect 7930 518 7982 570
rect 7994 518 8046 570
rect 8058 518 8110 570
rect 11504 518 11556 570
rect 11568 518 11620 570
rect 11632 518 11684 570
rect 11696 518 11748 570
rect 11760 518 11812 570
rect 15206 518 15258 570
rect 15270 518 15322 570
rect 15334 518 15386 570
rect 15398 518 15450 570
rect 15462 518 15514 570
<< metal2 >>
rect 1214 15600 1270 16000
rect 3146 15600 3202 16000
rect 5078 15600 5134 16000
rect 7010 15722 7066 16000
rect 8942 15722 8998 16000
rect 7010 15694 7144 15722
rect 7010 15600 7066 15694
rect 1228 14958 1256 15600
rect 2249 15260 2557 15269
rect 2249 15258 2255 15260
rect 2311 15258 2335 15260
rect 2391 15258 2415 15260
rect 2471 15258 2495 15260
rect 2551 15258 2557 15260
rect 2311 15206 2313 15258
rect 2493 15206 2495 15258
rect 2249 15204 2255 15206
rect 2311 15204 2335 15206
rect 2391 15204 2415 15206
rect 2471 15204 2495 15206
rect 2551 15204 2557 15206
rect 2249 15195 2557 15204
rect 3160 14958 3188 15600
rect 5092 14958 5120 15600
rect 5951 15260 6259 15269
rect 5951 15258 5957 15260
rect 6013 15258 6037 15260
rect 6093 15258 6117 15260
rect 6173 15258 6197 15260
rect 6253 15258 6259 15260
rect 6013 15206 6015 15258
rect 6195 15206 6197 15258
rect 5951 15204 5957 15206
rect 6013 15204 6037 15206
rect 6093 15204 6117 15206
rect 6173 15204 6197 15206
rect 6253 15204 6259 15206
rect 5951 15195 6259 15204
rect 7116 14958 7144 15694
rect 8772 15694 8998 15722
rect 8772 14958 8800 15694
rect 8942 15600 8998 15694
rect 10874 15722 10930 16000
rect 10874 15694 11008 15722
rect 10874 15600 10930 15694
rect 9653 15260 9961 15269
rect 9653 15258 9659 15260
rect 9715 15258 9739 15260
rect 9795 15258 9819 15260
rect 9875 15258 9899 15260
rect 9955 15258 9961 15260
rect 9715 15206 9717 15258
rect 9897 15206 9899 15258
rect 9653 15204 9659 15206
rect 9715 15204 9739 15206
rect 9795 15204 9819 15206
rect 9875 15204 9899 15206
rect 9955 15204 9961 15206
rect 9653 15195 9961 15204
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 1216 14952 1268 14958
rect 1216 14894 1268 14900
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 4528 14884 4580 14890
rect 4528 14826 4580 14832
rect 5632 14884 5684 14890
rect 5632 14826 5684 14832
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 1504 14618 1532 14758
rect 3988 14618 4016 14758
rect 4100 14716 4408 14725
rect 4100 14714 4106 14716
rect 4162 14714 4186 14716
rect 4242 14714 4266 14716
rect 4322 14714 4346 14716
rect 4402 14714 4408 14716
rect 4162 14662 4164 14714
rect 4344 14662 4346 14714
rect 4100 14660 4106 14662
rect 4162 14660 4186 14662
rect 4242 14660 4266 14662
rect 4322 14660 4346 14662
rect 4402 14660 4408 14662
rect 4100 14651 4408 14660
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 2249 14172 2557 14181
rect 2249 14170 2255 14172
rect 2311 14170 2335 14172
rect 2391 14170 2415 14172
rect 2471 14170 2495 14172
rect 2551 14170 2557 14172
rect 2311 14118 2313 14170
rect 2493 14118 2495 14170
rect 2249 14116 2255 14118
rect 2311 14116 2335 14118
rect 2391 14116 2415 14118
rect 2471 14116 2495 14118
rect 2551 14116 2557 14118
rect 2249 14107 2557 14116
rect 3988 14074 4016 14554
rect 4448 14482 4476 14758
rect 4540 14550 4568 14826
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4528 14544 4580 14550
rect 4528 14486 4580 14492
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 4540 14074 4568 14282
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4100 13628 4408 13637
rect 4100 13626 4106 13628
rect 4162 13626 4186 13628
rect 4242 13626 4266 13628
rect 4322 13626 4346 13628
rect 4402 13626 4408 13628
rect 4162 13574 4164 13626
rect 4344 13574 4346 13626
rect 4100 13572 4106 13574
rect 4162 13572 4186 13574
rect 4242 13572 4266 13574
rect 4322 13572 4346 13574
rect 4402 13572 4408 13574
rect 4100 13563 4408 13572
rect 4632 13530 4660 14418
rect 4724 13870 4752 14758
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5172 14340 5224 14346
rect 5172 14282 5224 14288
rect 5184 13938 5212 14282
rect 5368 14226 5396 14418
rect 5276 14198 5396 14226
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 5276 13870 5304 14198
rect 5460 14074 5488 14418
rect 5644 14346 5672 14826
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 5632 14340 5684 14346
rect 5632 14282 5684 14288
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 2249 13084 2557 13093
rect 2249 13082 2255 13084
rect 2311 13082 2335 13084
rect 2391 13082 2415 13084
rect 2471 13082 2495 13084
rect 2551 13082 2557 13084
rect 2311 13030 2313 13082
rect 2493 13030 2495 13082
rect 2249 13028 2255 13030
rect 2311 13028 2335 13030
rect 2391 13028 2415 13030
rect 2471 13028 2495 13030
rect 2551 13028 2557 13030
rect 2249 13019 2557 13028
rect 4724 12986 4752 13806
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 4804 13252 4856 13258
rect 4804 13194 4856 13200
rect 4816 12986 4844 13194
rect 5184 12986 5212 13262
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4100 12540 4408 12549
rect 4100 12538 4106 12540
rect 4162 12538 4186 12540
rect 4242 12538 4266 12540
rect 4322 12538 4346 12540
rect 4402 12538 4408 12540
rect 4162 12486 4164 12538
rect 4344 12486 4346 12538
rect 4100 12484 4106 12486
rect 4162 12484 4186 12486
rect 4242 12484 4266 12486
rect 4322 12484 4346 12486
rect 4402 12484 4408 12486
rect 4100 12475 4408 12484
rect 4724 12442 4752 12922
rect 5276 12782 5304 13806
rect 5828 13734 5856 14214
rect 5951 14172 6259 14181
rect 5951 14170 5957 14172
rect 6013 14170 6037 14172
rect 6093 14170 6117 14172
rect 6173 14170 6197 14172
rect 6253 14170 6259 14172
rect 6013 14118 6015 14170
rect 6195 14118 6197 14170
rect 5951 14116 5957 14118
rect 6013 14116 6037 14118
rect 6093 14116 6117 14118
rect 6173 14116 6197 14118
rect 6253 14116 6259 14118
rect 5951 14107 6259 14116
rect 6288 14074 6316 14758
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6380 13870 6408 14350
rect 6564 14346 6592 14894
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 7802 14716 8110 14725
rect 7802 14714 7808 14716
rect 7864 14714 7888 14716
rect 7944 14714 7968 14716
rect 8024 14714 8048 14716
rect 8104 14714 8110 14716
rect 7864 14662 7866 14714
rect 8046 14662 8048 14714
rect 7802 14660 7808 14662
rect 7864 14660 7888 14662
rect 7944 14660 7968 14662
rect 8024 14660 8048 14662
rect 8104 14660 8110 14662
rect 7802 14651 8110 14660
rect 8772 14618 8800 14758
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 6552 14340 6604 14346
rect 6552 14282 6604 14288
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 5368 13394 5396 13670
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5368 12442 5396 13330
rect 5951 13084 6259 13093
rect 5951 13082 5957 13084
rect 6013 13082 6037 13084
rect 6093 13082 6117 13084
rect 6173 13082 6197 13084
rect 6253 13082 6259 13084
rect 6013 13030 6015 13082
rect 6195 13030 6197 13082
rect 5951 13028 5957 13030
rect 6013 13028 6037 13030
rect 6093 13028 6117 13030
rect 6173 13028 6197 13030
rect 6253 13028 6259 13030
rect 5951 13019 6259 13028
rect 6748 12986 6776 13670
rect 7116 13190 7144 14418
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 5356 12436 5408 12442
rect 5920 12434 5948 12718
rect 6748 12646 6776 12922
rect 7116 12850 7144 13126
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7012 12776 7064 12782
rect 7208 12730 7236 14010
rect 7392 14006 7420 14214
rect 7576 14074 7604 14418
rect 8404 14074 8432 14418
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 8680 13870 8708 14554
rect 9324 14278 9352 14758
rect 9416 14550 9444 15098
rect 10980 15026 11008 15694
rect 12806 15600 12862 16000
rect 14738 15600 14794 16000
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 12820 14958 12848 15600
rect 13355 15260 13663 15269
rect 13355 15258 13361 15260
rect 13417 15258 13441 15260
rect 13497 15258 13521 15260
rect 13577 15258 13601 15260
rect 13657 15258 13663 15260
rect 13417 15206 13419 15258
rect 13599 15206 13601 15258
rect 13355 15204 13361 15206
rect 13417 15204 13441 15206
rect 13497 15204 13521 15206
rect 13577 15204 13601 15206
rect 13657 15204 13663 15206
rect 13355 15195 13663 15204
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 9692 14618 9720 14894
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 10336 14618 10364 14758
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 9404 14544 9456 14550
rect 9404 14486 9456 14492
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 7802 13628 8110 13637
rect 7802 13626 7808 13628
rect 7864 13626 7888 13628
rect 7944 13626 7968 13628
rect 8024 13626 8048 13628
rect 8104 13626 8110 13628
rect 7864 13574 7866 13626
rect 8046 13574 8048 13626
rect 7802 13572 7808 13574
rect 7864 13572 7888 13574
rect 7944 13572 7968 13574
rect 8024 13572 8048 13574
rect 8104 13572 8110 13574
rect 7802 13563 8110 13572
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7012 12718 7064 12724
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 5356 12378 5408 12384
rect 5828 12406 5948 12434
rect 5828 12102 5856 12406
rect 7024 12102 7052 12718
rect 7116 12702 7236 12730
rect 7116 12442 7144 12702
rect 7392 12458 7420 13330
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7852 12714 7880 13126
rect 7840 12708 7892 12714
rect 7840 12650 7892 12656
rect 7802 12540 8110 12549
rect 7802 12538 7808 12540
rect 7864 12538 7888 12540
rect 7944 12538 7968 12540
rect 8024 12538 8048 12540
rect 8104 12538 8110 12540
rect 7864 12486 7866 12538
rect 8046 12486 8048 12538
rect 7802 12484 7808 12486
rect 7864 12484 7888 12486
rect 7944 12484 7968 12486
rect 8024 12484 8048 12486
rect 8104 12484 8110 12486
rect 7802 12475 8110 12484
rect 7208 12442 7420 12458
rect 8220 12442 8248 13806
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7196 12436 7420 12442
rect 7248 12430 7420 12436
rect 8208 12436 8260 12442
rect 7196 12378 7248 12384
rect 8208 12378 8260 12384
rect 8404 12306 8432 12582
rect 9324 12306 9352 14214
rect 9416 14074 9444 14486
rect 10428 14278 10456 14758
rect 11504 14716 11812 14725
rect 11504 14714 11510 14716
rect 11566 14714 11590 14716
rect 11646 14714 11670 14716
rect 11726 14714 11750 14716
rect 11806 14714 11812 14716
rect 11566 14662 11568 14714
rect 11748 14662 11750 14714
rect 11504 14660 11510 14662
rect 11566 14660 11590 14662
rect 11646 14660 11670 14662
rect 11726 14660 11750 14662
rect 11806 14660 11812 14662
rect 11504 14651 11812 14660
rect 11900 14498 11928 14758
rect 11808 14470 11928 14498
rect 11808 14414 11836 14470
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9508 13938 9536 14214
rect 9653 14172 9961 14181
rect 9653 14170 9659 14172
rect 9715 14170 9739 14172
rect 9795 14170 9819 14172
rect 9875 14170 9899 14172
rect 9955 14170 9961 14172
rect 9715 14118 9717 14170
rect 9897 14118 9899 14170
rect 9653 14116 9659 14118
rect 9715 14116 9739 14118
rect 9795 14116 9819 14118
rect 9875 14116 9899 14118
rect 9955 14116 9961 14118
rect 9653 14107 9961 14116
rect 10428 14074 10456 14214
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 9784 13394 9812 13738
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10060 13462 10088 13670
rect 11256 13530 11284 13738
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10888 13258 10916 13330
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 9653 13084 9961 13093
rect 9653 13082 9659 13084
rect 9715 13082 9739 13084
rect 9795 13082 9819 13084
rect 9875 13082 9899 13084
rect 9955 13082 9961 13084
rect 9715 13030 9717 13082
rect 9897 13030 9899 13082
rect 9653 13028 9659 13030
rect 9715 13028 9739 13030
rect 9795 13028 9819 13030
rect 9875 13028 9899 13030
rect 9955 13028 9961 13030
rect 9653 13019 9961 13028
rect 10888 12986 10916 13194
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 11348 12782 11376 14350
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 9404 12708 9456 12714
rect 9404 12650 9456 12656
rect 9416 12442 9444 12650
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 2249 11996 2557 12005
rect 2249 11994 2255 11996
rect 2311 11994 2335 11996
rect 2391 11994 2415 11996
rect 2471 11994 2495 11996
rect 2551 11994 2557 11996
rect 2311 11942 2313 11994
rect 2493 11942 2495 11994
rect 2249 11940 2255 11942
rect 2311 11940 2335 11942
rect 2391 11940 2415 11942
rect 2471 11940 2495 11942
rect 2551 11940 2557 11942
rect 2249 11931 2557 11940
rect 5951 11996 6259 12005
rect 5951 11994 5957 11996
rect 6013 11994 6037 11996
rect 6093 11994 6117 11996
rect 6173 11994 6197 11996
rect 6253 11994 6259 11996
rect 6013 11942 6015 11994
rect 6195 11942 6197 11994
rect 5951 11940 5957 11942
rect 6013 11940 6037 11942
rect 6093 11940 6117 11942
rect 6173 11940 6197 11942
rect 6253 11940 6259 11942
rect 5951 11931 6259 11940
rect 9653 11996 9961 12005
rect 9653 11994 9659 11996
rect 9715 11994 9739 11996
rect 9795 11994 9819 11996
rect 9875 11994 9899 11996
rect 9955 11994 9961 11996
rect 9715 11942 9717 11994
rect 9897 11942 9899 11994
rect 9653 11940 9659 11942
rect 9715 11940 9739 11942
rect 9795 11940 9819 11942
rect 9875 11940 9899 11942
rect 9955 11940 9961 11942
rect 9653 11931 9961 11940
rect 4100 11452 4408 11461
rect 4100 11450 4106 11452
rect 4162 11450 4186 11452
rect 4242 11450 4266 11452
rect 4322 11450 4346 11452
rect 4402 11450 4408 11452
rect 4162 11398 4164 11450
rect 4344 11398 4346 11450
rect 4100 11396 4106 11398
rect 4162 11396 4186 11398
rect 4242 11396 4266 11398
rect 4322 11396 4346 11398
rect 4402 11396 4408 11398
rect 4100 11387 4408 11396
rect 7802 11452 8110 11461
rect 7802 11450 7808 11452
rect 7864 11450 7888 11452
rect 7944 11450 7968 11452
rect 8024 11450 8048 11452
rect 8104 11450 8110 11452
rect 7864 11398 7866 11450
rect 8046 11398 8048 11450
rect 7802 11396 7808 11398
rect 7864 11396 7888 11398
rect 7944 11396 7968 11398
rect 8024 11396 8048 11398
rect 8104 11396 8110 11398
rect 7802 11387 8110 11396
rect 2249 10908 2557 10917
rect 2249 10906 2255 10908
rect 2311 10906 2335 10908
rect 2391 10906 2415 10908
rect 2471 10906 2495 10908
rect 2551 10906 2557 10908
rect 2311 10854 2313 10906
rect 2493 10854 2495 10906
rect 2249 10852 2255 10854
rect 2311 10852 2335 10854
rect 2391 10852 2415 10854
rect 2471 10852 2495 10854
rect 2551 10852 2557 10854
rect 2249 10843 2557 10852
rect 5951 10908 6259 10917
rect 5951 10906 5957 10908
rect 6013 10906 6037 10908
rect 6093 10906 6117 10908
rect 6173 10906 6197 10908
rect 6253 10906 6259 10908
rect 6013 10854 6015 10906
rect 6195 10854 6197 10906
rect 5951 10852 5957 10854
rect 6013 10852 6037 10854
rect 6093 10852 6117 10854
rect 6173 10852 6197 10854
rect 6253 10852 6259 10854
rect 5951 10843 6259 10852
rect 9653 10908 9961 10917
rect 9653 10906 9659 10908
rect 9715 10906 9739 10908
rect 9795 10906 9819 10908
rect 9875 10906 9899 10908
rect 9955 10906 9961 10908
rect 9715 10854 9717 10906
rect 9897 10854 9899 10906
rect 9653 10852 9659 10854
rect 9715 10852 9739 10854
rect 9795 10852 9819 10854
rect 9875 10852 9899 10854
rect 9955 10852 9961 10854
rect 9653 10843 9961 10852
rect 4100 10364 4408 10373
rect 4100 10362 4106 10364
rect 4162 10362 4186 10364
rect 4242 10362 4266 10364
rect 4322 10362 4346 10364
rect 4402 10362 4408 10364
rect 4162 10310 4164 10362
rect 4344 10310 4346 10362
rect 4100 10308 4106 10310
rect 4162 10308 4186 10310
rect 4242 10308 4266 10310
rect 4322 10308 4346 10310
rect 4402 10308 4408 10310
rect 4100 10299 4408 10308
rect 7802 10364 8110 10373
rect 7802 10362 7808 10364
rect 7864 10362 7888 10364
rect 7944 10362 7968 10364
rect 8024 10362 8048 10364
rect 8104 10362 8110 10364
rect 7864 10310 7866 10362
rect 8046 10310 8048 10362
rect 7802 10308 7808 10310
rect 7864 10308 7888 10310
rect 7944 10308 7968 10310
rect 8024 10308 8048 10310
rect 8104 10308 8110 10310
rect 7802 10299 8110 10308
rect 2249 9820 2557 9829
rect 2249 9818 2255 9820
rect 2311 9818 2335 9820
rect 2391 9818 2415 9820
rect 2471 9818 2495 9820
rect 2551 9818 2557 9820
rect 2311 9766 2313 9818
rect 2493 9766 2495 9818
rect 2249 9764 2255 9766
rect 2311 9764 2335 9766
rect 2391 9764 2415 9766
rect 2471 9764 2495 9766
rect 2551 9764 2557 9766
rect 2249 9755 2557 9764
rect 5951 9820 6259 9829
rect 5951 9818 5957 9820
rect 6013 9818 6037 9820
rect 6093 9818 6117 9820
rect 6173 9818 6197 9820
rect 6253 9818 6259 9820
rect 6013 9766 6015 9818
rect 6195 9766 6197 9818
rect 5951 9764 5957 9766
rect 6013 9764 6037 9766
rect 6093 9764 6117 9766
rect 6173 9764 6197 9766
rect 6253 9764 6259 9766
rect 5951 9755 6259 9764
rect 9653 9820 9961 9829
rect 9653 9818 9659 9820
rect 9715 9818 9739 9820
rect 9795 9818 9819 9820
rect 9875 9818 9899 9820
rect 9955 9818 9961 9820
rect 9715 9766 9717 9818
rect 9897 9766 9899 9818
rect 9653 9764 9659 9766
rect 9715 9764 9739 9766
rect 9795 9764 9819 9766
rect 9875 9764 9899 9766
rect 9955 9764 9961 9766
rect 9653 9755 9961 9764
rect 4100 9276 4408 9285
rect 4100 9274 4106 9276
rect 4162 9274 4186 9276
rect 4242 9274 4266 9276
rect 4322 9274 4346 9276
rect 4402 9274 4408 9276
rect 4162 9222 4164 9274
rect 4344 9222 4346 9274
rect 4100 9220 4106 9222
rect 4162 9220 4186 9222
rect 4242 9220 4266 9222
rect 4322 9220 4346 9222
rect 4402 9220 4408 9222
rect 4100 9211 4408 9220
rect 7802 9276 8110 9285
rect 7802 9274 7808 9276
rect 7864 9274 7888 9276
rect 7944 9274 7968 9276
rect 8024 9274 8048 9276
rect 8104 9274 8110 9276
rect 7864 9222 7866 9274
rect 8046 9222 8048 9274
rect 7802 9220 7808 9222
rect 7864 9220 7888 9222
rect 7944 9220 7968 9222
rect 8024 9220 8048 9222
rect 8104 9220 8110 9222
rect 7802 9211 8110 9220
rect 2249 8732 2557 8741
rect 2249 8730 2255 8732
rect 2311 8730 2335 8732
rect 2391 8730 2415 8732
rect 2471 8730 2495 8732
rect 2551 8730 2557 8732
rect 2311 8678 2313 8730
rect 2493 8678 2495 8730
rect 2249 8676 2255 8678
rect 2311 8676 2335 8678
rect 2391 8676 2415 8678
rect 2471 8676 2495 8678
rect 2551 8676 2557 8678
rect 2249 8667 2557 8676
rect 5951 8732 6259 8741
rect 5951 8730 5957 8732
rect 6013 8730 6037 8732
rect 6093 8730 6117 8732
rect 6173 8730 6197 8732
rect 6253 8730 6259 8732
rect 6013 8678 6015 8730
rect 6195 8678 6197 8730
rect 5951 8676 5957 8678
rect 6013 8676 6037 8678
rect 6093 8676 6117 8678
rect 6173 8676 6197 8678
rect 6253 8676 6259 8678
rect 5951 8667 6259 8676
rect 9653 8732 9961 8741
rect 9653 8730 9659 8732
rect 9715 8730 9739 8732
rect 9795 8730 9819 8732
rect 9875 8730 9899 8732
rect 9955 8730 9961 8732
rect 9715 8678 9717 8730
rect 9897 8678 9899 8730
rect 9653 8676 9659 8678
rect 9715 8676 9739 8678
rect 9795 8676 9819 8678
rect 9875 8676 9899 8678
rect 9955 8676 9961 8678
rect 9653 8667 9961 8676
rect 4100 8188 4408 8197
rect 4100 8186 4106 8188
rect 4162 8186 4186 8188
rect 4242 8186 4266 8188
rect 4322 8186 4346 8188
rect 4402 8186 4408 8188
rect 4162 8134 4164 8186
rect 4344 8134 4346 8186
rect 4100 8132 4106 8134
rect 4162 8132 4186 8134
rect 4242 8132 4266 8134
rect 4322 8132 4346 8134
rect 4402 8132 4408 8134
rect 4100 8123 4408 8132
rect 7802 8188 8110 8197
rect 7802 8186 7808 8188
rect 7864 8186 7888 8188
rect 7944 8186 7968 8188
rect 8024 8186 8048 8188
rect 8104 8186 8110 8188
rect 7864 8134 7866 8186
rect 8046 8134 8048 8186
rect 7802 8132 7808 8134
rect 7864 8132 7888 8134
rect 7944 8132 7968 8134
rect 8024 8132 8048 8134
rect 8104 8132 8110 8134
rect 7802 8123 8110 8132
rect 2249 7644 2557 7653
rect 2249 7642 2255 7644
rect 2311 7642 2335 7644
rect 2391 7642 2415 7644
rect 2471 7642 2495 7644
rect 2551 7642 2557 7644
rect 2311 7590 2313 7642
rect 2493 7590 2495 7642
rect 2249 7588 2255 7590
rect 2311 7588 2335 7590
rect 2391 7588 2415 7590
rect 2471 7588 2495 7590
rect 2551 7588 2557 7590
rect 2249 7579 2557 7588
rect 5951 7644 6259 7653
rect 5951 7642 5957 7644
rect 6013 7642 6037 7644
rect 6093 7642 6117 7644
rect 6173 7642 6197 7644
rect 6253 7642 6259 7644
rect 6013 7590 6015 7642
rect 6195 7590 6197 7642
rect 5951 7588 5957 7590
rect 6013 7588 6037 7590
rect 6093 7588 6117 7590
rect 6173 7588 6197 7590
rect 6253 7588 6259 7590
rect 5951 7579 6259 7588
rect 9653 7644 9961 7653
rect 9653 7642 9659 7644
rect 9715 7642 9739 7644
rect 9795 7642 9819 7644
rect 9875 7642 9899 7644
rect 9955 7642 9961 7644
rect 9715 7590 9717 7642
rect 9897 7590 9899 7642
rect 9653 7588 9659 7590
rect 9715 7588 9739 7590
rect 9795 7588 9819 7590
rect 9875 7588 9899 7590
rect 9955 7588 9961 7590
rect 9653 7579 9961 7588
rect 4100 7100 4408 7109
rect 4100 7098 4106 7100
rect 4162 7098 4186 7100
rect 4242 7098 4266 7100
rect 4322 7098 4346 7100
rect 4402 7098 4408 7100
rect 4162 7046 4164 7098
rect 4344 7046 4346 7098
rect 4100 7044 4106 7046
rect 4162 7044 4186 7046
rect 4242 7044 4266 7046
rect 4322 7044 4346 7046
rect 4402 7044 4408 7046
rect 4100 7035 4408 7044
rect 7802 7100 8110 7109
rect 7802 7098 7808 7100
rect 7864 7098 7888 7100
rect 7944 7098 7968 7100
rect 8024 7098 8048 7100
rect 8104 7098 8110 7100
rect 7864 7046 7866 7098
rect 8046 7046 8048 7098
rect 7802 7044 7808 7046
rect 7864 7044 7888 7046
rect 7944 7044 7968 7046
rect 8024 7044 8048 7046
rect 8104 7044 8110 7046
rect 7802 7035 8110 7044
rect 11440 6914 11468 14010
rect 11992 13938 12020 14826
rect 12452 14074 12480 14894
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13096 14482 13124 14758
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12452 13938 12480 14010
rect 13280 13938 13308 14214
rect 13355 14172 13663 14181
rect 13355 14170 13361 14172
rect 13417 14170 13441 14172
rect 13497 14170 13521 14172
rect 13577 14170 13601 14172
rect 13657 14170 13663 14172
rect 13417 14118 13419 14170
rect 13599 14118 13601 14170
rect 13355 14116 13361 14118
rect 13417 14116 13441 14118
rect 13497 14116 13521 14118
rect 13577 14116 13601 14118
rect 13657 14116 13663 14118
rect 13355 14107 13663 14116
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11504 13628 11812 13637
rect 11504 13626 11510 13628
rect 11566 13626 11590 13628
rect 11646 13626 11670 13628
rect 11726 13626 11750 13628
rect 11806 13626 11812 13628
rect 11566 13574 11568 13626
rect 11748 13574 11750 13626
rect 11504 13572 11510 13574
rect 11566 13572 11590 13574
rect 11646 13572 11670 13574
rect 11726 13572 11750 13574
rect 11806 13572 11812 13574
rect 11504 13563 11812 13572
rect 11900 13326 11928 13806
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 12268 13530 12296 13670
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12268 12782 12296 13126
rect 12256 12776 12308 12782
rect 12256 12718 12308 12724
rect 13280 12714 13308 13670
rect 13355 13084 13663 13093
rect 13355 13082 13361 13084
rect 13417 13082 13441 13084
rect 13497 13082 13521 13084
rect 13577 13082 13601 13084
rect 13657 13082 13663 13084
rect 13417 13030 13419 13082
rect 13599 13030 13601 13082
rect 13355 13028 13361 13030
rect 13417 13028 13441 13030
rect 13497 13028 13521 13030
rect 13577 13028 13601 13030
rect 13657 13028 13663 13030
rect 13355 13019 13663 13028
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 11504 12540 11812 12549
rect 11504 12538 11510 12540
rect 11566 12538 11590 12540
rect 11646 12538 11670 12540
rect 11726 12538 11750 12540
rect 11806 12538 11812 12540
rect 11566 12486 11568 12538
rect 11748 12486 11750 12538
rect 11504 12484 11510 12486
rect 11566 12484 11590 12486
rect 11646 12484 11670 12486
rect 11726 12484 11750 12486
rect 11806 12484 11812 12486
rect 11504 12475 11812 12484
rect 13832 12306 13860 14554
rect 14752 14006 14780 15600
rect 15206 14716 15514 14725
rect 15206 14714 15212 14716
rect 15268 14714 15292 14716
rect 15348 14714 15372 14716
rect 15428 14714 15452 14716
rect 15508 14714 15514 14716
rect 15268 14662 15270 14714
rect 15450 14662 15452 14714
rect 15206 14660 15212 14662
rect 15268 14660 15292 14662
rect 15348 14660 15372 14662
rect 15428 14660 15452 14662
rect 15508 14660 15514 14662
rect 15206 14651 15514 14660
rect 14740 14000 14792 14006
rect 14740 13942 14792 13948
rect 15206 13628 15514 13637
rect 15206 13626 15212 13628
rect 15268 13626 15292 13628
rect 15348 13626 15372 13628
rect 15428 13626 15452 13628
rect 15508 13626 15514 13628
rect 15268 13574 15270 13626
rect 15450 13574 15452 13626
rect 15206 13572 15212 13574
rect 15268 13572 15292 13574
rect 15348 13572 15372 13574
rect 15428 13572 15452 13574
rect 15508 13572 15514 13574
rect 15206 13563 15514 13572
rect 15206 12540 15514 12549
rect 15206 12538 15212 12540
rect 15268 12538 15292 12540
rect 15348 12538 15372 12540
rect 15428 12538 15452 12540
rect 15508 12538 15514 12540
rect 15268 12486 15270 12538
rect 15450 12486 15452 12538
rect 15206 12484 15212 12486
rect 15268 12484 15292 12486
rect 15348 12484 15372 12486
rect 15428 12484 15452 12486
rect 15508 12484 15514 12486
rect 15206 12475 15514 12484
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 13355 11996 13663 12005
rect 13355 11994 13361 11996
rect 13417 11994 13441 11996
rect 13497 11994 13521 11996
rect 13577 11994 13601 11996
rect 13657 11994 13663 11996
rect 13417 11942 13419 11994
rect 13599 11942 13601 11994
rect 13355 11940 13361 11942
rect 13417 11940 13441 11942
rect 13497 11940 13521 11942
rect 13577 11940 13601 11942
rect 13657 11940 13663 11942
rect 13355 11931 13663 11940
rect 14752 11801 14780 12038
rect 14738 11792 14794 11801
rect 14738 11727 14794 11736
rect 11504 11452 11812 11461
rect 11504 11450 11510 11452
rect 11566 11450 11590 11452
rect 11646 11450 11670 11452
rect 11726 11450 11750 11452
rect 11806 11450 11812 11452
rect 11566 11398 11568 11450
rect 11748 11398 11750 11450
rect 11504 11396 11510 11398
rect 11566 11396 11590 11398
rect 11646 11396 11670 11398
rect 11726 11396 11750 11398
rect 11806 11396 11812 11398
rect 11504 11387 11812 11396
rect 15206 11452 15514 11461
rect 15206 11450 15212 11452
rect 15268 11450 15292 11452
rect 15348 11450 15372 11452
rect 15428 11450 15452 11452
rect 15508 11450 15514 11452
rect 15268 11398 15270 11450
rect 15450 11398 15452 11450
rect 15206 11396 15212 11398
rect 15268 11396 15292 11398
rect 15348 11396 15372 11398
rect 15428 11396 15452 11398
rect 15508 11396 15514 11398
rect 15206 11387 15514 11396
rect 13355 10908 13663 10917
rect 13355 10906 13361 10908
rect 13417 10906 13441 10908
rect 13497 10906 13521 10908
rect 13577 10906 13601 10908
rect 13657 10906 13663 10908
rect 13417 10854 13419 10906
rect 13599 10854 13601 10906
rect 13355 10852 13361 10854
rect 13417 10852 13441 10854
rect 13497 10852 13521 10854
rect 13577 10852 13601 10854
rect 13657 10852 13663 10854
rect 13355 10843 13663 10852
rect 11504 10364 11812 10373
rect 11504 10362 11510 10364
rect 11566 10362 11590 10364
rect 11646 10362 11670 10364
rect 11726 10362 11750 10364
rect 11806 10362 11812 10364
rect 11566 10310 11568 10362
rect 11748 10310 11750 10362
rect 11504 10308 11510 10310
rect 11566 10308 11590 10310
rect 11646 10308 11670 10310
rect 11726 10308 11750 10310
rect 11806 10308 11812 10310
rect 11504 10299 11812 10308
rect 15206 10364 15514 10373
rect 15206 10362 15212 10364
rect 15268 10362 15292 10364
rect 15348 10362 15372 10364
rect 15428 10362 15452 10364
rect 15508 10362 15514 10364
rect 15268 10310 15270 10362
rect 15450 10310 15452 10362
rect 15206 10308 15212 10310
rect 15268 10308 15292 10310
rect 15348 10308 15372 10310
rect 15428 10308 15452 10310
rect 15508 10308 15514 10310
rect 15206 10299 15514 10308
rect 13355 9820 13663 9829
rect 13355 9818 13361 9820
rect 13417 9818 13441 9820
rect 13497 9818 13521 9820
rect 13577 9818 13601 9820
rect 13657 9818 13663 9820
rect 13417 9766 13419 9818
rect 13599 9766 13601 9818
rect 13355 9764 13361 9766
rect 13417 9764 13441 9766
rect 13497 9764 13521 9766
rect 13577 9764 13601 9766
rect 13657 9764 13663 9766
rect 13355 9755 13663 9764
rect 11504 9276 11812 9285
rect 11504 9274 11510 9276
rect 11566 9274 11590 9276
rect 11646 9274 11670 9276
rect 11726 9274 11750 9276
rect 11806 9274 11812 9276
rect 11566 9222 11568 9274
rect 11748 9222 11750 9274
rect 11504 9220 11510 9222
rect 11566 9220 11590 9222
rect 11646 9220 11670 9222
rect 11726 9220 11750 9222
rect 11806 9220 11812 9222
rect 11504 9211 11812 9220
rect 15206 9276 15514 9285
rect 15206 9274 15212 9276
rect 15268 9274 15292 9276
rect 15348 9274 15372 9276
rect 15428 9274 15452 9276
rect 15508 9274 15514 9276
rect 15268 9222 15270 9274
rect 15450 9222 15452 9274
rect 15206 9220 15212 9222
rect 15268 9220 15292 9222
rect 15348 9220 15372 9222
rect 15428 9220 15452 9222
rect 15508 9220 15514 9222
rect 15206 9211 15514 9220
rect 13355 8732 13663 8741
rect 13355 8730 13361 8732
rect 13417 8730 13441 8732
rect 13497 8730 13521 8732
rect 13577 8730 13601 8732
rect 13657 8730 13663 8732
rect 13417 8678 13419 8730
rect 13599 8678 13601 8730
rect 13355 8676 13361 8678
rect 13417 8676 13441 8678
rect 13497 8676 13521 8678
rect 13577 8676 13601 8678
rect 13657 8676 13663 8678
rect 13355 8667 13663 8676
rect 11504 8188 11812 8197
rect 11504 8186 11510 8188
rect 11566 8186 11590 8188
rect 11646 8186 11670 8188
rect 11726 8186 11750 8188
rect 11806 8186 11812 8188
rect 11566 8134 11568 8186
rect 11748 8134 11750 8186
rect 11504 8132 11510 8134
rect 11566 8132 11590 8134
rect 11646 8132 11670 8134
rect 11726 8132 11750 8134
rect 11806 8132 11812 8134
rect 11504 8123 11812 8132
rect 15206 8188 15514 8197
rect 15206 8186 15212 8188
rect 15268 8186 15292 8188
rect 15348 8186 15372 8188
rect 15428 8186 15452 8188
rect 15508 8186 15514 8188
rect 15268 8134 15270 8186
rect 15450 8134 15452 8186
rect 15206 8132 15212 8134
rect 15268 8132 15292 8134
rect 15348 8132 15372 8134
rect 15428 8132 15452 8134
rect 15508 8132 15514 8134
rect 15206 8123 15514 8132
rect 13355 7644 13663 7653
rect 13355 7642 13361 7644
rect 13417 7642 13441 7644
rect 13497 7642 13521 7644
rect 13577 7642 13601 7644
rect 13657 7642 13663 7644
rect 13417 7590 13419 7642
rect 13599 7590 13601 7642
rect 13355 7588 13361 7590
rect 13417 7588 13441 7590
rect 13497 7588 13521 7590
rect 13577 7588 13601 7590
rect 13657 7588 13663 7590
rect 13355 7579 13663 7588
rect 11504 7100 11812 7109
rect 11504 7098 11510 7100
rect 11566 7098 11590 7100
rect 11646 7098 11670 7100
rect 11726 7098 11750 7100
rect 11806 7098 11812 7100
rect 11566 7046 11568 7098
rect 11748 7046 11750 7098
rect 11504 7044 11510 7046
rect 11566 7044 11590 7046
rect 11646 7044 11670 7046
rect 11726 7044 11750 7046
rect 11806 7044 11812 7046
rect 11504 7035 11812 7044
rect 15206 7100 15514 7109
rect 15206 7098 15212 7100
rect 15268 7098 15292 7100
rect 15348 7098 15372 7100
rect 15428 7098 15452 7100
rect 15508 7098 15514 7100
rect 15268 7046 15270 7098
rect 15450 7046 15452 7098
rect 15206 7044 15212 7046
rect 15268 7044 15292 7046
rect 15348 7044 15372 7046
rect 15428 7044 15452 7046
rect 15508 7044 15514 7046
rect 15206 7035 15514 7044
rect 11348 6886 11468 6914
rect 2249 6556 2557 6565
rect 2249 6554 2255 6556
rect 2311 6554 2335 6556
rect 2391 6554 2415 6556
rect 2471 6554 2495 6556
rect 2551 6554 2557 6556
rect 2311 6502 2313 6554
rect 2493 6502 2495 6554
rect 2249 6500 2255 6502
rect 2311 6500 2335 6502
rect 2391 6500 2415 6502
rect 2471 6500 2495 6502
rect 2551 6500 2557 6502
rect 2249 6491 2557 6500
rect 5951 6556 6259 6565
rect 5951 6554 5957 6556
rect 6013 6554 6037 6556
rect 6093 6554 6117 6556
rect 6173 6554 6197 6556
rect 6253 6554 6259 6556
rect 6013 6502 6015 6554
rect 6195 6502 6197 6554
rect 5951 6500 5957 6502
rect 6013 6500 6037 6502
rect 6093 6500 6117 6502
rect 6173 6500 6197 6502
rect 6253 6500 6259 6502
rect 5951 6491 6259 6500
rect 9653 6556 9961 6565
rect 9653 6554 9659 6556
rect 9715 6554 9739 6556
rect 9795 6554 9819 6556
rect 9875 6554 9899 6556
rect 9955 6554 9961 6556
rect 9715 6502 9717 6554
rect 9897 6502 9899 6554
rect 9653 6500 9659 6502
rect 9715 6500 9739 6502
rect 9795 6500 9819 6502
rect 9875 6500 9899 6502
rect 9955 6500 9961 6502
rect 9653 6491 9961 6500
rect 4100 6012 4408 6021
rect 4100 6010 4106 6012
rect 4162 6010 4186 6012
rect 4242 6010 4266 6012
rect 4322 6010 4346 6012
rect 4402 6010 4408 6012
rect 4162 5958 4164 6010
rect 4344 5958 4346 6010
rect 4100 5956 4106 5958
rect 4162 5956 4186 5958
rect 4242 5956 4266 5958
rect 4322 5956 4346 5958
rect 4402 5956 4408 5958
rect 4100 5947 4408 5956
rect 7802 6012 8110 6021
rect 7802 6010 7808 6012
rect 7864 6010 7888 6012
rect 7944 6010 7968 6012
rect 8024 6010 8048 6012
rect 8104 6010 8110 6012
rect 7864 5958 7866 6010
rect 8046 5958 8048 6010
rect 7802 5956 7808 5958
rect 7864 5956 7888 5958
rect 7944 5956 7968 5958
rect 8024 5956 8048 5958
rect 8104 5956 8110 5958
rect 7802 5947 8110 5956
rect 2249 5468 2557 5477
rect 2249 5466 2255 5468
rect 2311 5466 2335 5468
rect 2391 5466 2415 5468
rect 2471 5466 2495 5468
rect 2551 5466 2557 5468
rect 2311 5414 2313 5466
rect 2493 5414 2495 5466
rect 2249 5412 2255 5414
rect 2311 5412 2335 5414
rect 2391 5412 2415 5414
rect 2471 5412 2495 5414
rect 2551 5412 2557 5414
rect 2249 5403 2557 5412
rect 5951 5468 6259 5477
rect 5951 5466 5957 5468
rect 6013 5466 6037 5468
rect 6093 5466 6117 5468
rect 6173 5466 6197 5468
rect 6253 5466 6259 5468
rect 6013 5414 6015 5466
rect 6195 5414 6197 5466
rect 5951 5412 5957 5414
rect 6013 5412 6037 5414
rect 6093 5412 6117 5414
rect 6173 5412 6197 5414
rect 6253 5412 6259 5414
rect 5951 5403 6259 5412
rect 9653 5468 9961 5477
rect 9653 5466 9659 5468
rect 9715 5466 9739 5468
rect 9795 5466 9819 5468
rect 9875 5466 9899 5468
rect 9955 5466 9961 5468
rect 9715 5414 9717 5466
rect 9897 5414 9899 5466
rect 9653 5412 9659 5414
rect 9715 5412 9739 5414
rect 9795 5412 9819 5414
rect 9875 5412 9899 5414
rect 9955 5412 9961 5414
rect 9653 5403 9961 5412
rect 4100 4924 4408 4933
rect 4100 4922 4106 4924
rect 4162 4922 4186 4924
rect 4242 4922 4266 4924
rect 4322 4922 4346 4924
rect 4402 4922 4408 4924
rect 4162 4870 4164 4922
rect 4344 4870 4346 4922
rect 4100 4868 4106 4870
rect 4162 4868 4186 4870
rect 4242 4868 4266 4870
rect 4322 4868 4346 4870
rect 4402 4868 4408 4870
rect 4100 4859 4408 4868
rect 7802 4924 8110 4933
rect 7802 4922 7808 4924
rect 7864 4922 7888 4924
rect 7944 4922 7968 4924
rect 8024 4922 8048 4924
rect 8104 4922 8110 4924
rect 7864 4870 7866 4922
rect 8046 4870 8048 4922
rect 7802 4868 7808 4870
rect 7864 4868 7888 4870
rect 7944 4868 7968 4870
rect 8024 4868 8048 4870
rect 8104 4868 8110 4870
rect 7802 4859 8110 4868
rect 11348 4758 11376 6886
rect 13355 6556 13663 6565
rect 13355 6554 13361 6556
rect 13417 6554 13441 6556
rect 13497 6554 13521 6556
rect 13577 6554 13601 6556
rect 13657 6554 13663 6556
rect 13417 6502 13419 6554
rect 13599 6502 13601 6554
rect 13355 6500 13361 6502
rect 13417 6500 13441 6502
rect 13497 6500 13521 6502
rect 13577 6500 13601 6502
rect 13657 6500 13663 6502
rect 13355 6491 13663 6500
rect 11504 6012 11812 6021
rect 11504 6010 11510 6012
rect 11566 6010 11590 6012
rect 11646 6010 11670 6012
rect 11726 6010 11750 6012
rect 11806 6010 11812 6012
rect 11566 5958 11568 6010
rect 11748 5958 11750 6010
rect 11504 5956 11510 5958
rect 11566 5956 11590 5958
rect 11646 5956 11670 5958
rect 11726 5956 11750 5958
rect 11806 5956 11812 5958
rect 11504 5947 11812 5956
rect 15206 6012 15514 6021
rect 15206 6010 15212 6012
rect 15268 6010 15292 6012
rect 15348 6010 15372 6012
rect 15428 6010 15452 6012
rect 15508 6010 15514 6012
rect 15268 5958 15270 6010
rect 15450 5958 15452 6010
rect 15206 5956 15212 5958
rect 15268 5956 15292 5958
rect 15348 5956 15372 5958
rect 15428 5956 15452 5958
rect 15508 5956 15514 5958
rect 15206 5947 15514 5956
rect 13355 5468 13663 5477
rect 13355 5466 13361 5468
rect 13417 5466 13441 5468
rect 13497 5466 13521 5468
rect 13577 5466 13601 5468
rect 13657 5466 13663 5468
rect 13417 5414 13419 5466
rect 13599 5414 13601 5466
rect 13355 5412 13361 5414
rect 13417 5412 13441 5414
rect 13497 5412 13521 5414
rect 13577 5412 13601 5414
rect 13657 5412 13663 5414
rect 13355 5403 13663 5412
rect 11504 4924 11812 4933
rect 11504 4922 11510 4924
rect 11566 4922 11590 4924
rect 11646 4922 11670 4924
rect 11726 4922 11750 4924
rect 11806 4922 11812 4924
rect 11566 4870 11568 4922
rect 11748 4870 11750 4922
rect 11504 4868 11510 4870
rect 11566 4868 11590 4870
rect 11646 4868 11670 4870
rect 11726 4868 11750 4870
rect 11806 4868 11812 4870
rect 11504 4859 11812 4868
rect 15206 4924 15514 4933
rect 15206 4922 15212 4924
rect 15268 4922 15292 4924
rect 15348 4922 15372 4924
rect 15428 4922 15452 4924
rect 15508 4922 15514 4924
rect 15268 4870 15270 4922
rect 15450 4870 15452 4922
rect 15206 4868 15212 4870
rect 15268 4868 15292 4870
rect 15348 4868 15372 4870
rect 15428 4868 15452 4870
rect 15508 4868 15514 4870
rect 15206 4859 15514 4868
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 2249 4380 2557 4389
rect 2249 4378 2255 4380
rect 2311 4378 2335 4380
rect 2391 4378 2415 4380
rect 2471 4378 2495 4380
rect 2551 4378 2557 4380
rect 2311 4326 2313 4378
rect 2493 4326 2495 4378
rect 2249 4324 2255 4326
rect 2311 4324 2335 4326
rect 2391 4324 2415 4326
rect 2471 4324 2495 4326
rect 2551 4324 2557 4326
rect 2249 4315 2557 4324
rect 5951 4380 6259 4389
rect 5951 4378 5957 4380
rect 6013 4378 6037 4380
rect 6093 4378 6117 4380
rect 6173 4378 6197 4380
rect 6253 4378 6259 4380
rect 6013 4326 6015 4378
rect 6195 4326 6197 4378
rect 5951 4324 5957 4326
rect 6013 4324 6037 4326
rect 6093 4324 6117 4326
rect 6173 4324 6197 4326
rect 6253 4324 6259 4326
rect 5951 4315 6259 4324
rect 9653 4380 9961 4389
rect 9653 4378 9659 4380
rect 9715 4378 9739 4380
rect 9795 4378 9819 4380
rect 9875 4378 9899 4380
rect 9955 4378 9961 4380
rect 9715 4326 9717 4378
rect 9897 4326 9899 4378
rect 9653 4324 9659 4326
rect 9715 4324 9739 4326
rect 9795 4324 9819 4326
rect 9875 4324 9899 4326
rect 9955 4324 9961 4326
rect 9653 4315 9961 4324
rect 11256 4185 11284 4422
rect 13355 4380 13663 4389
rect 13355 4378 13361 4380
rect 13417 4378 13441 4380
rect 13497 4378 13521 4380
rect 13577 4378 13601 4380
rect 13657 4378 13663 4380
rect 13417 4326 13419 4378
rect 13599 4326 13601 4378
rect 13355 4324 13361 4326
rect 13417 4324 13441 4326
rect 13497 4324 13521 4326
rect 13577 4324 13601 4326
rect 13657 4324 13663 4326
rect 13355 4315 13663 4324
rect 11242 4176 11298 4185
rect 11242 4111 11298 4120
rect 4100 3836 4408 3845
rect 4100 3834 4106 3836
rect 4162 3834 4186 3836
rect 4242 3834 4266 3836
rect 4322 3834 4346 3836
rect 4402 3834 4408 3836
rect 4162 3782 4164 3834
rect 4344 3782 4346 3834
rect 4100 3780 4106 3782
rect 4162 3780 4186 3782
rect 4242 3780 4266 3782
rect 4322 3780 4346 3782
rect 4402 3780 4408 3782
rect 4100 3771 4408 3780
rect 7802 3836 8110 3845
rect 7802 3834 7808 3836
rect 7864 3834 7888 3836
rect 7944 3834 7968 3836
rect 8024 3834 8048 3836
rect 8104 3834 8110 3836
rect 7864 3782 7866 3834
rect 8046 3782 8048 3834
rect 7802 3780 7808 3782
rect 7864 3780 7888 3782
rect 7944 3780 7968 3782
rect 8024 3780 8048 3782
rect 8104 3780 8110 3782
rect 7802 3771 8110 3780
rect 11504 3836 11812 3845
rect 11504 3834 11510 3836
rect 11566 3834 11590 3836
rect 11646 3834 11670 3836
rect 11726 3834 11750 3836
rect 11806 3834 11812 3836
rect 11566 3782 11568 3834
rect 11748 3782 11750 3834
rect 11504 3780 11510 3782
rect 11566 3780 11590 3782
rect 11646 3780 11670 3782
rect 11726 3780 11750 3782
rect 11806 3780 11812 3782
rect 11504 3771 11812 3780
rect 15206 3836 15514 3845
rect 15206 3834 15212 3836
rect 15268 3834 15292 3836
rect 15348 3834 15372 3836
rect 15428 3834 15452 3836
rect 15508 3834 15514 3836
rect 15268 3782 15270 3834
rect 15450 3782 15452 3834
rect 15206 3780 15212 3782
rect 15268 3780 15292 3782
rect 15348 3780 15372 3782
rect 15428 3780 15452 3782
rect 15508 3780 15514 3782
rect 15206 3771 15514 3780
rect 2249 3292 2557 3301
rect 2249 3290 2255 3292
rect 2311 3290 2335 3292
rect 2391 3290 2415 3292
rect 2471 3290 2495 3292
rect 2551 3290 2557 3292
rect 2311 3238 2313 3290
rect 2493 3238 2495 3290
rect 2249 3236 2255 3238
rect 2311 3236 2335 3238
rect 2391 3236 2415 3238
rect 2471 3236 2495 3238
rect 2551 3236 2557 3238
rect 2249 3227 2557 3236
rect 5951 3292 6259 3301
rect 5951 3290 5957 3292
rect 6013 3290 6037 3292
rect 6093 3290 6117 3292
rect 6173 3290 6197 3292
rect 6253 3290 6259 3292
rect 6013 3238 6015 3290
rect 6195 3238 6197 3290
rect 5951 3236 5957 3238
rect 6013 3236 6037 3238
rect 6093 3236 6117 3238
rect 6173 3236 6197 3238
rect 6253 3236 6259 3238
rect 5951 3227 6259 3236
rect 9653 3292 9961 3301
rect 9653 3290 9659 3292
rect 9715 3290 9739 3292
rect 9795 3290 9819 3292
rect 9875 3290 9899 3292
rect 9955 3290 9961 3292
rect 9715 3238 9717 3290
rect 9897 3238 9899 3290
rect 9653 3236 9659 3238
rect 9715 3236 9739 3238
rect 9795 3236 9819 3238
rect 9875 3236 9899 3238
rect 9955 3236 9961 3238
rect 9653 3227 9961 3236
rect 13355 3292 13663 3301
rect 13355 3290 13361 3292
rect 13417 3290 13441 3292
rect 13497 3290 13521 3292
rect 13577 3290 13601 3292
rect 13657 3290 13663 3292
rect 13417 3238 13419 3290
rect 13599 3238 13601 3290
rect 13355 3236 13361 3238
rect 13417 3236 13441 3238
rect 13497 3236 13521 3238
rect 13577 3236 13601 3238
rect 13657 3236 13663 3238
rect 13355 3227 13663 3236
rect 4100 2748 4408 2757
rect 4100 2746 4106 2748
rect 4162 2746 4186 2748
rect 4242 2746 4266 2748
rect 4322 2746 4346 2748
rect 4402 2746 4408 2748
rect 4162 2694 4164 2746
rect 4344 2694 4346 2746
rect 4100 2692 4106 2694
rect 4162 2692 4186 2694
rect 4242 2692 4266 2694
rect 4322 2692 4346 2694
rect 4402 2692 4408 2694
rect 4100 2683 4408 2692
rect 7802 2748 8110 2757
rect 7802 2746 7808 2748
rect 7864 2746 7888 2748
rect 7944 2746 7968 2748
rect 8024 2746 8048 2748
rect 8104 2746 8110 2748
rect 7864 2694 7866 2746
rect 8046 2694 8048 2746
rect 7802 2692 7808 2694
rect 7864 2692 7888 2694
rect 7944 2692 7968 2694
rect 8024 2692 8048 2694
rect 8104 2692 8110 2694
rect 7802 2683 8110 2692
rect 11504 2748 11812 2757
rect 11504 2746 11510 2748
rect 11566 2746 11590 2748
rect 11646 2746 11670 2748
rect 11726 2746 11750 2748
rect 11806 2746 11812 2748
rect 11566 2694 11568 2746
rect 11748 2694 11750 2746
rect 11504 2692 11510 2694
rect 11566 2692 11590 2694
rect 11646 2692 11670 2694
rect 11726 2692 11750 2694
rect 11806 2692 11812 2694
rect 11504 2683 11812 2692
rect 15206 2748 15514 2757
rect 15206 2746 15212 2748
rect 15268 2746 15292 2748
rect 15348 2746 15372 2748
rect 15428 2746 15452 2748
rect 15508 2746 15514 2748
rect 15268 2694 15270 2746
rect 15450 2694 15452 2746
rect 15206 2692 15212 2694
rect 15268 2692 15292 2694
rect 15348 2692 15372 2694
rect 15428 2692 15452 2694
rect 15508 2692 15514 2694
rect 15206 2683 15514 2692
rect 2249 2204 2557 2213
rect 2249 2202 2255 2204
rect 2311 2202 2335 2204
rect 2391 2202 2415 2204
rect 2471 2202 2495 2204
rect 2551 2202 2557 2204
rect 2311 2150 2313 2202
rect 2493 2150 2495 2202
rect 2249 2148 2255 2150
rect 2311 2148 2335 2150
rect 2391 2148 2415 2150
rect 2471 2148 2495 2150
rect 2551 2148 2557 2150
rect 2249 2139 2557 2148
rect 5951 2204 6259 2213
rect 5951 2202 5957 2204
rect 6013 2202 6037 2204
rect 6093 2202 6117 2204
rect 6173 2202 6197 2204
rect 6253 2202 6259 2204
rect 6013 2150 6015 2202
rect 6195 2150 6197 2202
rect 5951 2148 5957 2150
rect 6013 2148 6037 2150
rect 6093 2148 6117 2150
rect 6173 2148 6197 2150
rect 6253 2148 6259 2150
rect 5951 2139 6259 2148
rect 9653 2204 9961 2213
rect 9653 2202 9659 2204
rect 9715 2202 9739 2204
rect 9795 2202 9819 2204
rect 9875 2202 9899 2204
rect 9955 2202 9961 2204
rect 9715 2150 9717 2202
rect 9897 2150 9899 2202
rect 9653 2148 9659 2150
rect 9715 2148 9739 2150
rect 9795 2148 9819 2150
rect 9875 2148 9899 2150
rect 9955 2148 9961 2150
rect 9653 2139 9961 2148
rect 13355 2204 13663 2213
rect 13355 2202 13361 2204
rect 13417 2202 13441 2204
rect 13497 2202 13521 2204
rect 13577 2202 13601 2204
rect 13657 2202 13663 2204
rect 13417 2150 13419 2202
rect 13599 2150 13601 2202
rect 13355 2148 13361 2150
rect 13417 2148 13441 2150
rect 13497 2148 13521 2150
rect 13577 2148 13601 2150
rect 13657 2148 13663 2150
rect 13355 2139 13663 2148
rect 4100 1660 4408 1669
rect 4100 1658 4106 1660
rect 4162 1658 4186 1660
rect 4242 1658 4266 1660
rect 4322 1658 4346 1660
rect 4402 1658 4408 1660
rect 4162 1606 4164 1658
rect 4344 1606 4346 1658
rect 4100 1604 4106 1606
rect 4162 1604 4186 1606
rect 4242 1604 4266 1606
rect 4322 1604 4346 1606
rect 4402 1604 4408 1606
rect 4100 1595 4408 1604
rect 7802 1660 8110 1669
rect 7802 1658 7808 1660
rect 7864 1658 7888 1660
rect 7944 1658 7968 1660
rect 8024 1658 8048 1660
rect 8104 1658 8110 1660
rect 7864 1606 7866 1658
rect 8046 1606 8048 1658
rect 7802 1604 7808 1606
rect 7864 1604 7888 1606
rect 7944 1604 7968 1606
rect 8024 1604 8048 1606
rect 8104 1604 8110 1606
rect 7802 1595 8110 1604
rect 11504 1660 11812 1669
rect 11504 1658 11510 1660
rect 11566 1658 11590 1660
rect 11646 1658 11670 1660
rect 11726 1658 11750 1660
rect 11806 1658 11812 1660
rect 11566 1606 11568 1658
rect 11748 1606 11750 1658
rect 11504 1604 11510 1606
rect 11566 1604 11590 1606
rect 11646 1604 11670 1606
rect 11726 1604 11750 1606
rect 11806 1604 11812 1606
rect 11504 1595 11812 1604
rect 15206 1660 15514 1669
rect 15206 1658 15212 1660
rect 15268 1658 15292 1660
rect 15348 1658 15372 1660
rect 15428 1658 15452 1660
rect 15508 1658 15514 1660
rect 15268 1606 15270 1658
rect 15450 1606 15452 1658
rect 15206 1604 15212 1606
rect 15268 1604 15292 1606
rect 15348 1604 15372 1606
rect 15428 1604 15452 1606
rect 15508 1604 15514 1606
rect 15206 1595 15514 1604
rect 2249 1116 2557 1125
rect 2249 1114 2255 1116
rect 2311 1114 2335 1116
rect 2391 1114 2415 1116
rect 2471 1114 2495 1116
rect 2551 1114 2557 1116
rect 2311 1062 2313 1114
rect 2493 1062 2495 1114
rect 2249 1060 2255 1062
rect 2311 1060 2335 1062
rect 2391 1060 2415 1062
rect 2471 1060 2495 1062
rect 2551 1060 2557 1062
rect 2249 1051 2557 1060
rect 5951 1116 6259 1125
rect 5951 1114 5957 1116
rect 6013 1114 6037 1116
rect 6093 1114 6117 1116
rect 6173 1114 6197 1116
rect 6253 1114 6259 1116
rect 6013 1062 6015 1114
rect 6195 1062 6197 1114
rect 5951 1060 5957 1062
rect 6013 1060 6037 1062
rect 6093 1060 6117 1062
rect 6173 1060 6197 1062
rect 6253 1060 6259 1062
rect 5951 1051 6259 1060
rect 9653 1116 9961 1125
rect 9653 1114 9659 1116
rect 9715 1114 9739 1116
rect 9795 1114 9819 1116
rect 9875 1114 9899 1116
rect 9955 1114 9961 1116
rect 9715 1062 9717 1114
rect 9897 1062 9899 1114
rect 9653 1060 9659 1062
rect 9715 1060 9739 1062
rect 9795 1060 9819 1062
rect 9875 1060 9899 1062
rect 9955 1060 9961 1062
rect 9653 1051 9961 1060
rect 13355 1116 13663 1125
rect 13355 1114 13361 1116
rect 13417 1114 13441 1116
rect 13497 1114 13521 1116
rect 13577 1114 13601 1116
rect 13657 1114 13663 1116
rect 13417 1062 13419 1114
rect 13599 1062 13601 1114
rect 13355 1060 13361 1062
rect 13417 1060 13441 1062
rect 13497 1060 13521 1062
rect 13577 1060 13601 1062
rect 13657 1060 13663 1062
rect 13355 1051 13663 1060
rect 4100 572 4408 581
rect 4100 570 4106 572
rect 4162 570 4186 572
rect 4242 570 4266 572
rect 4322 570 4346 572
rect 4402 570 4408 572
rect 4162 518 4164 570
rect 4344 518 4346 570
rect 4100 516 4106 518
rect 4162 516 4186 518
rect 4242 516 4266 518
rect 4322 516 4346 518
rect 4402 516 4408 518
rect 4100 507 4408 516
rect 7802 572 8110 581
rect 7802 570 7808 572
rect 7864 570 7888 572
rect 7944 570 7968 572
rect 8024 570 8048 572
rect 8104 570 8110 572
rect 7864 518 7866 570
rect 8046 518 8048 570
rect 7802 516 7808 518
rect 7864 516 7888 518
rect 7944 516 7968 518
rect 8024 516 8048 518
rect 8104 516 8110 518
rect 7802 507 8110 516
rect 11504 572 11812 581
rect 11504 570 11510 572
rect 11566 570 11590 572
rect 11646 570 11670 572
rect 11726 570 11750 572
rect 11806 570 11812 572
rect 11566 518 11568 570
rect 11748 518 11750 570
rect 11504 516 11510 518
rect 11566 516 11590 518
rect 11646 516 11670 518
rect 11726 516 11750 518
rect 11806 516 11812 518
rect 11504 507 11812 516
rect 15206 572 15514 581
rect 15206 570 15212 572
rect 15268 570 15292 572
rect 15348 570 15372 572
rect 15428 570 15452 572
rect 15508 570 15514 572
rect 15268 518 15270 570
rect 15450 518 15452 570
rect 15206 516 15212 518
rect 15268 516 15292 518
rect 15348 516 15372 518
rect 15428 516 15452 518
rect 15508 516 15514 518
rect 15206 507 15514 516
<< via2 >>
rect 2255 15258 2311 15260
rect 2335 15258 2391 15260
rect 2415 15258 2471 15260
rect 2495 15258 2551 15260
rect 2255 15206 2301 15258
rect 2301 15206 2311 15258
rect 2335 15206 2365 15258
rect 2365 15206 2377 15258
rect 2377 15206 2391 15258
rect 2415 15206 2429 15258
rect 2429 15206 2441 15258
rect 2441 15206 2471 15258
rect 2495 15206 2505 15258
rect 2505 15206 2551 15258
rect 2255 15204 2311 15206
rect 2335 15204 2391 15206
rect 2415 15204 2471 15206
rect 2495 15204 2551 15206
rect 5957 15258 6013 15260
rect 6037 15258 6093 15260
rect 6117 15258 6173 15260
rect 6197 15258 6253 15260
rect 5957 15206 6003 15258
rect 6003 15206 6013 15258
rect 6037 15206 6067 15258
rect 6067 15206 6079 15258
rect 6079 15206 6093 15258
rect 6117 15206 6131 15258
rect 6131 15206 6143 15258
rect 6143 15206 6173 15258
rect 6197 15206 6207 15258
rect 6207 15206 6253 15258
rect 5957 15204 6013 15206
rect 6037 15204 6093 15206
rect 6117 15204 6173 15206
rect 6197 15204 6253 15206
rect 9659 15258 9715 15260
rect 9739 15258 9795 15260
rect 9819 15258 9875 15260
rect 9899 15258 9955 15260
rect 9659 15206 9705 15258
rect 9705 15206 9715 15258
rect 9739 15206 9769 15258
rect 9769 15206 9781 15258
rect 9781 15206 9795 15258
rect 9819 15206 9833 15258
rect 9833 15206 9845 15258
rect 9845 15206 9875 15258
rect 9899 15206 9909 15258
rect 9909 15206 9955 15258
rect 9659 15204 9715 15206
rect 9739 15204 9795 15206
rect 9819 15204 9875 15206
rect 9899 15204 9955 15206
rect 4106 14714 4162 14716
rect 4186 14714 4242 14716
rect 4266 14714 4322 14716
rect 4346 14714 4402 14716
rect 4106 14662 4152 14714
rect 4152 14662 4162 14714
rect 4186 14662 4216 14714
rect 4216 14662 4228 14714
rect 4228 14662 4242 14714
rect 4266 14662 4280 14714
rect 4280 14662 4292 14714
rect 4292 14662 4322 14714
rect 4346 14662 4356 14714
rect 4356 14662 4402 14714
rect 4106 14660 4162 14662
rect 4186 14660 4242 14662
rect 4266 14660 4322 14662
rect 4346 14660 4402 14662
rect 2255 14170 2311 14172
rect 2335 14170 2391 14172
rect 2415 14170 2471 14172
rect 2495 14170 2551 14172
rect 2255 14118 2301 14170
rect 2301 14118 2311 14170
rect 2335 14118 2365 14170
rect 2365 14118 2377 14170
rect 2377 14118 2391 14170
rect 2415 14118 2429 14170
rect 2429 14118 2441 14170
rect 2441 14118 2471 14170
rect 2495 14118 2505 14170
rect 2505 14118 2551 14170
rect 2255 14116 2311 14118
rect 2335 14116 2391 14118
rect 2415 14116 2471 14118
rect 2495 14116 2551 14118
rect 4106 13626 4162 13628
rect 4186 13626 4242 13628
rect 4266 13626 4322 13628
rect 4346 13626 4402 13628
rect 4106 13574 4152 13626
rect 4152 13574 4162 13626
rect 4186 13574 4216 13626
rect 4216 13574 4228 13626
rect 4228 13574 4242 13626
rect 4266 13574 4280 13626
rect 4280 13574 4292 13626
rect 4292 13574 4322 13626
rect 4346 13574 4356 13626
rect 4356 13574 4402 13626
rect 4106 13572 4162 13574
rect 4186 13572 4242 13574
rect 4266 13572 4322 13574
rect 4346 13572 4402 13574
rect 2255 13082 2311 13084
rect 2335 13082 2391 13084
rect 2415 13082 2471 13084
rect 2495 13082 2551 13084
rect 2255 13030 2301 13082
rect 2301 13030 2311 13082
rect 2335 13030 2365 13082
rect 2365 13030 2377 13082
rect 2377 13030 2391 13082
rect 2415 13030 2429 13082
rect 2429 13030 2441 13082
rect 2441 13030 2471 13082
rect 2495 13030 2505 13082
rect 2505 13030 2551 13082
rect 2255 13028 2311 13030
rect 2335 13028 2391 13030
rect 2415 13028 2471 13030
rect 2495 13028 2551 13030
rect 4106 12538 4162 12540
rect 4186 12538 4242 12540
rect 4266 12538 4322 12540
rect 4346 12538 4402 12540
rect 4106 12486 4152 12538
rect 4152 12486 4162 12538
rect 4186 12486 4216 12538
rect 4216 12486 4228 12538
rect 4228 12486 4242 12538
rect 4266 12486 4280 12538
rect 4280 12486 4292 12538
rect 4292 12486 4322 12538
rect 4346 12486 4356 12538
rect 4356 12486 4402 12538
rect 4106 12484 4162 12486
rect 4186 12484 4242 12486
rect 4266 12484 4322 12486
rect 4346 12484 4402 12486
rect 5957 14170 6013 14172
rect 6037 14170 6093 14172
rect 6117 14170 6173 14172
rect 6197 14170 6253 14172
rect 5957 14118 6003 14170
rect 6003 14118 6013 14170
rect 6037 14118 6067 14170
rect 6067 14118 6079 14170
rect 6079 14118 6093 14170
rect 6117 14118 6131 14170
rect 6131 14118 6143 14170
rect 6143 14118 6173 14170
rect 6197 14118 6207 14170
rect 6207 14118 6253 14170
rect 5957 14116 6013 14118
rect 6037 14116 6093 14118
rect 6117 14116 6173 14118
rect 6197 14116 6253 14118
rect 7808 14714 7864 14716
rect 7888 14714 7944 14716
rect 7968 14714 8024 14716
rect 8048 14714 8104 14716
rect 7808 14662 7854 14714
rect 7854 14662 7864 14714
rect 7888 14662 7918 14714
rect 7918 14662 7930 14714
rect 7930 14662 7944 14714
rect 7968 14662 7982 14714
rect 7982 14662 7994 14714
rect 7994 14662 8024 14714
rect 8048 14662 8058 14714
rect 8058 14662 8104 14714
rect 7808 14660 7864 14662
rect 7888 14660 7944 14662
rect 7968 14660 8024 14662
rect 8048 14660 8104 14662
rect 5957 13082 6013 13084
rect 6037 13082 6093 13084
rect 6117 13082 6173 13084
rect 6197 13082 6253 13084
rect 5957 13030 6003 13082
rect 6003 13030 6013 13082
rect 6037 13030 6067 13082
rect 6067 13030 6079 13082
rect 6079 13030 6093 13082
rect 6117 13030 6131 13082
rect 6131 13030 6143 13082
rect 6143 13030 6173 13082
rect 6197 13030 6207 13082
rect 6207 13030 6253 13082
rect 5957 13028 6013 13030
rect 6037 13028 6093 13030
rect 6117 13028 6173 13030
rect 6197 13028 6253 13030
rect 13361 15258 13417 15260
rect 13441 15258 13497 15260
rect 13521 15258 13577 15260
rect 13601 15258 13657 15260
rect 13361 15206 13407 15258
rect 13407 15206 13417 15258
rect 13441 15206 13471 15258
rect 13471 15206 13483 15258
rect 13483 15206 13497 15258
rect 13521 15206 13535 15258
rect 13535 15206 13547 15258
rect 13547 15206 13577 15258
rect 13601 15206 13611 15258
rect 13611 15206 13657 15258
rect 13361 15204 13417 15206
rect 13441 15204 13497 15206
rect 13521 15204 13577 15206
rect 13601 15204 13657 15206
rect 7808 13626 7864 13628
rect 7888 13626 7944 13628
rect 7968 13626 8024 13628
rect 8048 13626 8104 13628
rect 7808 13574 7854 13626
rect 7854 13574 7864 13626
rect 7888 13574 7918 13626
rect 7918 13574 7930 13626
rect 7930 13574 7944 13626
rect 7968 13574 7982 13626
rect 7982 13574 7994 13626
rect 7994 13574 8024 13626
rect 8048 13574 8058 13626
rect 8058 13574 8104 13626
rect 7808 13572 7864 13574
rect 7888 13572 7944 13574
rect 7968 13572 8024 13574
rect 8048 13572 8104 13574
rect 7808 12538 7864 12540
rect 7888 12538 7944 12540
rect 7968 12538 8024 12540
rect 8048 12538 8104 12540
rect 7808 12486 7854 12538
rect 7854 12486 7864 12538
rect 7888 12486 7918 12538
rect 7918 12486 7930 12538
rect 7930 12486 7944 12538
rect 7968 12486 7982 12538
rect 7982 12486 7994 12538
rect 7994 12486 8024 12538
rect 8048 12486 8058 12538
rect 8058 12486 8104 12538
rect 7808 12484 7864 12486
rect 7888 12484 7944 12486
rect 7968 12484 8024 12486
rect 8048 12484 8104 12486
rect 11510 14714 11566 14716
rect 11590 14714 11646 14716
rect 11670 14714 11726 14716
rect 11750 14714 11806 14716
rect 11510 14662 11556 14714
rect 11556 14662 11566 14714
rect 11590 14662 11620 14714
rect 11620 14662 11632 14714
rect 11632 14662 11646 14714
rect 11670 14662 11684 14714
rect 11684 14662 11696 14714
rect 11696 14662 11726 14714
rect 11750 14662 11760 14714
rect 11760 14662 11806 14714
rect 11510 14660 11566 14662
rect 11590 14660 11646 14662
rect 11670 14660 11726 14662
rect 11750 14660 11806 14662
rect 9659 14170 9715 14172
rect 9739 14170 9795 14172
rect 9819 14170 9875 14172
rect 9899 14170 9955 14172
rect 9659 14118 9705 14170
rect 9705 14118 9715 14170
rect 9739 14118 9769 14170
rect 9769 14118 9781 14170
rect 9781 14118 9795 14170
rect 9819 14118 9833 14170
rect 9833 14118 9845 14170
rect 9845 14118 9875 14170
rect 9899 14118 9909 14170
rect 9909 14118 9955 14170
rect 9659 14116 9715 14118
rect 9739 14116 9795 14118
rect 9819 14116 9875 14118
rect 9899 14116 9955 14118
rect 9659 13082 9715 13084
rect 9739 13082 9795 13084
rect 9819 13082 9875 13084
rect 9899 13082 9955 13084
rect 9659 13030 9705 13082
rect 9705 13030 9715 13082
rect 9739 13030 9769 13082
rect 9769 13030 9781 13082
rect 9781 13030 9795 13082
rect 9819 13030 9833 13082
rect 9833 13030 9845 13082
rect 9845 13030 9875 13082
rect 9899 13030 9909 13082
rect 9909 13030 9955 13082
rect 9659 13028 9715 13030
rect 9739 13028 9795 13030
rect 9819 13028 9875 13030
rect 9899 13028 9955 13030
rect 2255 11994 2311 11996
rect 2335 11994 2391 11996
rect 2415 11994 2471 11996
rect 2495 11994 2551 11996
rect 2255 11942 2301 11994
rect 2301 11942 2311 11994
rect 2335 11942 2365 11994
rect 2365 11942 2377 11994
rect 2377 11942 2391 11994
rect 2415 11942 2429 11994
rect 2429 11942 2441 11994
rect 2441 11942 2471 11994
rect 2495 11942 2505 11994
rect 2505 11942 2551 11994
rect 2255 11940 2311 11942
rect 2335 11940 2391 11942
rect 2415 11940 2471 11942
rect 2495 11940 2551 11942
rect 5957 11994 6013 11996
rect 6037 11994 6093 11996
rect 6117 11994 6173 11996
rect 6197 11994 6253 11996
rect 5957 11942 6003 11994
rect 6003 11942 6013 11994
rect 6037 11942 6067 11994
rect 6067 11942 6079 11994
rect 6079 11942 6093 11994
rect 6117 11942 6131 11994
rect 6131 11942 6143 11994
rect 6143 11942 6173 11994
rect 6197 11942 6207 11994
rect 6207 11942 6253 11994
rect 5957 11940 6013 11942
rect 6037 11940 6093 11942
rect 6117 11940 6173 11942
rect 6197 11940 6253 11942
rect 9659 11994 9715 11996
rect 9739 11994 9795 11996
rect 9819 11994 9875 11996
rect 9899 11994 9955 11996
rect 9659 11942 9705 11994
rect 9705 11942 9715 11994
rect 9739 11942 9769 11994
rect 9769 11942 9781 11994
rect 9781 11942 9795 11994
rect 9819 11942 9833 11994
rect 9833 11942 9845 11994
rect 9845 11942 9875 11994
rect 9899 11942 9909 11994
rect 9909 11942 9955 11994
rect 9659 11940 9715 11942
rect 9739 11940 9795 11942
rect 9819 11940 9875 11942
rect 9899 11940 9955 11942
rect 4106 11450 4162 11452
rect 4186 11450 4242 11452
rect 4266 11450 4322 11452
rect 4346 11450 4402 11452
rect 4106 11398 4152 11450
rect 4152 11398 4162 11450
rect 4186 11398 4216 11450
rect 4216 11398 4228 11450
rect 4228 11398 4242 11450
rect 4266 11398 4280 11450
rect 4280 11398 4292 11450
rect 4292 11398 4322 11450
rect 4346 11398 4356 11450
rect 4356 11398 4402 11450
rect 4106 11396 4162 11398
rect 4186 11396 4242 11398
rect 4266 11396 4322 11398
rect 4346 11396 4402 11398
rect 7808 11450 7864 11452
rect 7888 11450 7944 11452
rect 7968 11450 8024 11452
rect 8048 11450 8104 11452
rect 7808 11398 7854 11450
rect 7854 11398 7864 11450
rect 7888 11398 7918 11450
rect 7918 11398 7930 11450
rect 7930 11398 7944 11450
rect 7968 11398 7982 11450
rect 7982 11398 7994 11450
rect 7994 11398 8024 11450
rect 8048 11398 8058 11450
rect 8058 11398 8104 11450
rect 7808 11396 7864 11398
rect 7888 11396 7944 11398
rect 7968 11396 8024 11398
rect 8048 11396 8104 11398
rect 2255 10906 2311 10908
rect 2335 10906 2391 10908
rect 2415 10906 2471 10908
rect 2495 10906 2551 10908
rect 2255 10854 2301 10906
rect 2301 10854 2311 10906
rect 2335 10854 2365 10906
rect 2365 10854 2377 10906
rect 2377 10854 2391 10906
rect 2415 10854 2429 10906
rect 2429 10854 2441 10906
rect 2441 10854 2471 10906
rect 2495 10854 2505 10906
rect 2505 10854 2551 10906
rect 2255 10852 2311 10854
rect 2335 10852 2391 10854
rect 2415 10852 2471 10854
rect 2495 10852 2551 10854
rect 5957 10906 6013 10908
rect 6037 10906 6093 10908
rect 6117 10906 6173 10908
rect 6197 10906 6253 10908
rect 5957 10854 6003 10906
rect 6003 10854 6013 10906
rect 6037 10854 6067 10906
rect 6067 10854 6079 10906
rect 6079 10854 6093 10906
rect 6117 10854 6131 10906
rect 6131 10854 6143 10906
rect 6143 10854 6173 10906
rect 6197 10854 6207 10906
rect 6207 10854 6253 10906
rect 5957 10852 6013 10854
rect 6037 10852 6093 10854
rect 6117 10852 6173 10854
rect 6197 10852 6253 10854
rect 9659 10906 9715 10908
rect 9739 10906 9795 10908
rect 9819 10906 9875 10908
rect 9899 10906 9955 10908
rect 9659 10854 9705 10906
rect 9705 10854 9715 10906
rect 9739 10854 9769 10906
rect 9769 10854 9781 10906
rect 9781 10854 9795 10906
rect 9819 10854 9833 10906
rect 9833 10854 9845 10906
rect 9845 10854 9875 10906
rect 9899 10854 9909 10906
rect 9909 10854 9955 10906
rect 9659 10852 9715 10854
rect 9739 10852 9795 10854
rect 9819 10852 9875 10854
rect 9899 10852 9955 10854
rect 4106 10362 4162 10364
rect 4186 10362 4242 10364
rect 4266 10362 4322 10364
rect 4346 10362 4402 10364
rect 4106 10310 4152 10362
rect 4152 10310 4162 10362
rect 4186 10310 4216 10362
rect 4216 10310 4228 10362
rect 4228 10310 4242 10362
rect 4266 10310 4280 10362
rect 4280 10310 4292 10362
rect 4292 10310 4322 10362
rect 4346 10310 4356 10362
rect 4356 10310 4402 10362
rect 4106 10308 4162 10310
rect 4186 10308 4242 10310
rect 4266 10308 4322 10310
rect 4346 10308 4402 10310
rect 7808 10362 7864 10364
rect 7888 10362 7944 10364
rect 7968 10362 8024 10364
rect 8048 10362 8104 10364
rect 7808 10310 7854 10362
rect 7854 10310 7864 10362
rect 7888 10310 7918 10362
rect 7918 10310 7930 10362
rect 7930 10310 7944 10362
rect 7968 10310 7982 10362
rect 7982 10310 7994 10362
rect 7994 10310 8024 10362
rect 8048 10310 8058 10362
rect 8058 10310 8104 10362
rect 7808 10308 7864 10310
rect 7888 10308 7944 10310
rect 7968 10308 8024 10310
rect 8048 10308 8104 10310
rect 2255 9818 2311 9820
rect 2335 9818 2391 9820
rect 2415 9818 2471 9820
rect 2495 9818 2551 9820
rect 2255 9766 2301 9818
rect 2301 9766 2311 9818
rect 2335 9766 2365 9818
rect 2365 9766 2377 9818
rect 2377 9766 2391 9818
rect 2415 9766 2429 9818
rect 2429 9766 2441 9818
rect 2441 9766 2471 9818
rect 2495 9766 2505 9818
rect 2505 9766 2551 9818
rect 2255 9764 2311 9766
rect 2335 9764 2391 9766
rect 2415 9764 2471 9766
rect 2495 9764 2551 9766
rect 5957 9818 6013 9820
rect 6037 9818 6093 9820
rect 6117 9818 6173 9820
rect 6197 9818 6253 9820
rect 5957 9766 6003 9818
rect 6003 9766 6013 9818
rect 6037 9766 6067 9818
rect 6067 9766 6079 9818
rect 6079 9766 6093 9818
rect 6117 9766 6131 9818
rect 6131 9766 6143 9818
rect 6143 9766 6173 9818
rect 6197 9766 6207 9818
rect 6207 9766 6253 9818
rect 5957 9764 6013 9766
rect 6037 9764 6093 9766
rect 6117 9764 6173 9766
rect 6197 9764 6253 9766
rect 9659 9818 9715 9820
rect 9739 9818 9795 9820
rect 9819 9818 9875 9820
rect 9899 9818 9955 9820
rect 9659 9766 9705 9818
rect 9705 9766 9715 9818
rect 9739 9766 9769 9818
rect 9769 9766 9781 9818
rect 9781 9766 9795 9818
rect 9819 9766 9833 9818
rect 9833 9766 9845 9818
rect 9845 9766 9875 9818
rect 9899 9766 9909 9818
rect 9909 9766 9955 9818
rect 9659 9764 9715 9766
rect 9739 9764 9795 9766
rect 9819 9764 9875 9766
rect 9899 9764 9955 9766
rect 4106 9274 4162 9276
rect 4186 9274 4242 9276
rect 4266 9274 4322 9276
rect 4346 9274 4402 9276
rect 4106 9222 4152 9274
rect 4152 9222 4162 9274
rect 4186 9222 4216 9274
rect 4216 9222 4228 9274
rect 4228 9222 4242 9274
rect 4266 9222 4280 9274
rect 4280 9222 4292 9274
rect 4292 9222 4322 9274
rect 4346 9222 4356 9274
rect 4356 9222 4402 9274
rect 4106 9220 4162 9222
rect 4186 9220 4242 9222
rect 4266 9220 4322 9222
rect 4346 9220 4402 9222
rect 7808 9274 7864 9276
rect 7888 9274 7944 9276
rect 7968 9274 8024 9276
rect 8048 9274 8104 9276
rect 7808 9222 7854 9274
rect 7854 9222 7864 9274
rect 7888 9222 7918 9274
rect 7918 9222 7930 9274
rect 7930 9222 7944 9274
rect 7968 9222 7982 9274
rect 7982 9222 7994 9274
rect 7994 9222 8024 9274
rect 8048 9222 8058 9274
rect 8058 9222 8104 9274
rect 7808 9220 7864 9222
rect 7888 9220 7944 9222
rect 7968 9220 8024 9222
rect 8048 9220 8104 9222
rect 2255 8730 2311 8732
rect 2335 8730 2391 8732
rect 2415 8730 2471 8732
rect 2495 8730 2551 8732
rect 2255 8678 2301 8730
rect 2301 8678 2311 8730
rect 2335 8678 2365 8730
rect 2365 8678 2377 8730
rect 2377 8678 2391 8730
rect 2415 8678 2429 8730
rect 2429 8678 2441 8730
rect 2441 8678 2471 8730
rect 2495 8678 2505 8730
rect 2505 8678 2551 8730
rect 2255 8676 2311 8678
rect 2335 8676 2391 8678
rect 2415 8676 2471 8678
rect 2495 8676 2551 8678
rect 5957 8730 6013 8732
rect 6037 8730 6093 8732
rect 6117 8730 6173 8732
rect 6197 8730 6253 8732
rect 5957 8678 6003 8730
rect 6003 8678 6013 8730
rect 6037 8678 6067 8730
rect 6067 8678 6079 8730
rect 6079 8678 6093 8730
rect 6117 8678 6131 8730
rect 6131 8678 6143 8730
rect 6143 8678 6173 8730
rect 6197 8678 6207 8730
rect 6207 8678 6253 8730
rect 5957 8676 6013 8678
rect 6037 8676 6093 8678
rect 6117 8676 6173 8678
rect 6197 8676 6253 8678
rect 9659 8730 9715 8732
rect 9739 8730 9795 8732
rect 9819 8730 9875 8732
rect 9899 8730 9955 8732
rect 9659 8678 9705 8730
rect 9705 8678 9715 8730
rect 9739 8678 9769 8730
rect 9769 8678 9781 8730
rect 9781 8678 9795 8730
rect 9819 8678 9833 8730
rect 9833 8678 9845 8730
rect 9845 8678 9875 8730
rect 9899 8678 9909 8730
rect 9909 8678 9955 8730
rect 9659 8676 9715 8678
rect 9739 8676 9795 8678
rect 9819 8676 9875 8678
rect 9899 8676 9955 8678
rect 4106 8186 4162 8188
rect 4186 8186 4242 8188
rect 4266 8186 4322 8188
rect 4346 8186 4402 8188
rect 4106 8134 4152 8186
rect 4152 8134 4162 8186
rect 4186 8134 4216 8186
rect 4216 8134 4228 8186
rect 4228 8134 4242 8186
rect 4266 8134 4280 8186
rect 4280 8134 4292 8186
rect 4292 8134 4322 8186
rect 4346 8134 4356 8186
rect 4356 8134 4402 8186
rect 4106 8132 4162 8134
rect 4186 8132 4242 8134
rect 4266 8132 4322 8134
rect 4346 8132 4402 8134
rect 7808 8186 7864 8188
rect 7888 8186 7944 8188
rect 7968 8186 8024 8188
rect 8048 8186 8104 8188
rect 7808 8134 7854 8186
rect 7854 8134 7864 8186
rect 7888 8134 7918 8186
rect 7918 8134 7930 8186
rect 7930 8134 7944 8186
rect 7968 8134 7982 8186
rect 7982 8134 7994 8186
rect 7994 8134 8024 8186
rect 8048 8134 8058 8186
rect 8058 8134 8104 8186
rect 7808 8132 7864 8134
rect 7888 8132 7944 8134
rect 7968 8132 8024 8134
rect 8048 8132 8104 8134
rect 2255 7642 2311 7644
rect 2335 7642 2391 7644
rect 2415 7642 2471 7644
rect 2495 7642 2551 7644
rect 2255 7590 2301 7642
rect 2301 7590 2311 7642
rect 2335 7590 2365 7642
rect 2365 7590 2377 7642
rect 2377 7590 2391 7642
rect 2415 7590 2429 7642
rect 2429 7590 2441 7642
rect 2441 7590 2471 7642
rect 2495 7590 2505 7642
rect 2505 7590 2551 7642
rect 2255 7588 2311 7590
rect 2335 7588 2391 7590
rect 2415 7588 2471 7590
rect 2495 7588 2551 7590
rect 5957 7642 6013 7644
rect 6037 7642 6093 7644
rect 6117 7642 6173 7644
rect 6197 7642 6253 7644
rect 5957 7590 6003 7642
rect 6003 7590 6013 7642
rect 6037 7590 6067 7642
rect 6067 7590 6079 7642
rect 6079 7590 6093 7642
rect 6117 7590 6131 7642
rect 6131 7590 6143 7642
rect 6143 7590 6173 7642
rect 6197 7590 6207 7642
rect 6207 7590 6253 7642
rect 5957 7588 6013 7590
rect 6037 7588 6093 7590
rect 6117 7588 6173 7590
rect 6197 7588 6253 7590
rect 9659 7642 9715 7644
rect 9739 7642 9795 7644
rect 9819 7642 9875 7644
rect 9899 7642 9955 7644
rect 9659 7590 9705 7642
rect 9705 7590 9715 7642
rect 9739 7590 9769 7642
rect 9769 7590 9781 7642
rect 9781 7590 9795 7642
rect 9819 7590 9833 7642
rect 9833 7590 9845 7642
rect 9845 7590 9875 7642
rect 9899 7590 9909 7642
rect 9909 7590 9955 7642
rect 9659 7588 9715 7590
rect 9739 7588 9795 7590
rect 9819 7588 9875 7590
rect 9899 7588 9955 7590
rect 4106 7098 4162 7100
rect 4186 7098 4242 7100
rect 4266 7098 4322 7100
rect 4346 7098 4402 7100
rect 4106 7046 4152 7098
rect 4152 7046 4162 7098
rect 4186 7046 4216 7098
rect 4216 7046 4228 7098
rect 4228 7046 4242 7098
rect 4266 7046 4280 7098
rect 4280 7046 4292 7098
rect 4292 7046 4322 7098
rect 4346 7046 4356 7098
rect 4356 7046 4402 7098
rect 4106 7044 4162 7046
rect 4186 7044 4242 7046
rect 4266 7044 4322 7046
rect 4346 7044 4402 7046
rect 7808 7098 7864 7100
rect 7888 7098 7944 7100
rect 7968 7098 8024 7100
rect 8048 7098 8104 7100
rect 7808 7046 7854 7098
rect 7854 7046 7864 7098
rect 7888 7046 7918 7098
rect 7918 7046 7930 7098
rect 7930 7046 7944 7098
rect 7968 7046 7982 7098
rect 7982 7046 7994 7098
rect 7994 7046 8024 7098
rect 8048 7046 8058 7098
rect 8058 7046 8104 7098
rect 7808 7044 7864 7046
rect 7888 7044 7944 7046
rect 7968 7044 8024 7046
rect 8048 7044 8104 7046
rect 13361 14170 13417 14172
rect 13441 14170 13497 14172
rect 13521 14170 13577 14172
rect 13601 14170 13657 14172
rect 13361 14118 13407 14170
rect 13407 14118 13417 14170
rect 13441 14118 13471 14170
rect 13471 14118 13483 14170
rect 13483 14118 13497 14170
rect 13521 14118 13535 14170
rect 13535 14118 13547 14170
rect 13547 14118 13577 14170
rect 13601 14118 13611 14170
rect 13611 14118 13657 14170
rect 13361 14116 13417 14118
rect 13441 14116 13497 14118
rect 13521 14116 13577 14118
rect 13601 14116 13657 14118
rect 11510 13626 11566 13628
rect 11590 13626 11646 13628
rect 11670 13626 11726 13628
rect 11750 13626 11806 13628
rect 11510 13574 11556 13626
rect 11556 13574 11566 13626
rect 11590 13574 11620 13626
rect 11620 13574 11632 13626
rect 11632 13574 11646 13626
rect 11670 13574 11684 13626
rect 11684 13574 11696 13626
rect 11696 13574 11726 13626
rect 11750 13574 11760 13626
rect 11760 13574 11806 13626
rect 11510 13572 11566 13574
rect 11590 13572 11646 13574
rect 11670 13572 11726 13574
rect 11750 13572 11806 13574
rect 13361 13082 13417 13084
rect 13441 13082 13497 13084
rect 13521 13082 13577 13084
rect 13601 13082 13657 13084
rect 13361 13030 13407 13082
rect 13407 13030 13417 13082
rect 13441 13030 13471 13082
rect 13471 13030 13483 13082
rect 13483 13030 13497 13082
rect 13521 13030 13535 13082
rect 13535 13030 13547 13082
rect 13547 13030 13577 13082
rect 13601 13030 13611 13082
rect 13611 13030 13657 13082
rect 13361 13028 13417 13030
rect 13441 13028 13497 13030
rect 13521 13028 13577 13030
rect 13601 13028 13657 13030
rect 11510 12538 11566 12540
rect 11590 12538 11646 12540
rect 11670 12538 11726 12540
rect 11750 12538 11806 12540
rect 11510 12486 11556 12538
rect 11556 12486 11566 12538
rect 11590 12486 11620 12538
rect 11620 12486 11632 12538
rect 11632 12486 11646 12538
rect 11670 12486 11684 12538
rect 11684 12486 11696 12538
rect 11696 12486 11726 12538
rect 11750 12486 11760 12538
rect 11760 12486 11806 12538
rect 11510 12484 11566 12486
rect 11590 12484 11646 12486
rect 11670 12484 11726 12486
rect 11750 12484 11806 12486
rect 15212 14714 15268 14716
rect 15292 14714 15348 14716
rect 15372 14714 15428 14716
rect 15452 14714 15508 14716
rect 15212 14662 15258 14714
rect 15258 14662 15268 14714
rect 15292 14662 15322 14714
rect 15322 14662 15334 14714
rect 15334 14662 15348 14714
rect 15372 14662 15386 14714
rect 15386 14662 15398 14714
rect 15398 14662 15428 14714
rect 15452 14662 15462 14714
rect 15462 14662 15508 14714
rect 15212 14660 15268 14662
rect 15292 14660 15348 14662
rect 15372 14660 15428 14662
rect 15452 14660 15508 14662
rect 15212 13626 15268 13628
rect 15292 13626 15348 13628
rect 15372 13626 15428 13628
rect 15452 13626 15508 13628
rect 15212 13574 15258 13626
rect 15258 13574 15268 13626
rect 15292 13574 15322 13626
rect 15322 13574 15334 13626
rect 15334 13574 15348 13626
rect 15372 13574 15386 13626
rect 15386 13574 15398 13626
rect 15398 13574 15428 13626
rect 15452 13574 15462 13626
rect 15462 13574 15508 13626
rect 15212 13572 15268 13574
rect 15292 13572 15348 13574
rect 15372 13572 15428 13574
rect 15452 13572 15508 13574
rect 15212 12538 15268 12540
rect 15292 12538 15348 12540
rect 15372 12538 15428 12540
rect 15452 12538 15508 12540
rect 15212 12486 15258 12538
rect 15258 12486 15268 12538
rect 15292 12486 15322 12538
rect 15322 12486 15334 12538
rect 15334 12486 15348 12538
rect 15372 12486 15386 12538
rect 15386 12486 15398 12538
rect 15398 12486 15428 12538
rect 15452 12486 15462 12538
rect 15462 12486 15508 12538
rect 15212 12484 15268 12486
rect 15292 12484 15348 12486
rect 15372 12484 15428 12486
rect 15452 12484 15508 12486
rect 13361 11994 13417 11996
rect 13441 11994 13497 11996
rect 13521 11994 13577 11996
rect 13601 11994 13657 11996
rect 13361 11942 13407 11994
rect 13407 11942 13417 11994
rect 13441 11942 13471 11994
rect 13471 11942 13483 11994
rect 13483 11942 13497 11994
rect 13521 11942 13535 11994
rect 13535 11942 13547 11994
rect 13547 11942 13577 11994
rect 13601 11942 13611 11994
rect 13611 11942 13657 11994
rect 13361 11940 13417 11942
rect 13441 11940 13497 11942
rect 13521 11940 13577 11942
rect 13601 11940 13657 11942
rect 14738 11736 14794 11792
rect 11510 11450 11566 11452
rect 11590 11450 11646 11452
rect 11670 11450 11726 11452
rect 11750 11450 11806 11452
rect 11510 11398 11556 11450
rect 11556 11398 11566 11450
rect 11590 11398 11620 11450
rect 11620 11398 11632 11450
rect 11632 11398 11646 11450
rect 11670 11398 11684 11450
rect 11684 11398 11696 11450
rect 11696 11398 11726 11450
rect 11750 11398 11760 11450
rect 11760 11398 11806 11450
rect 11510 11396 11566 11398
rect 11590 11396 11646 11398
rect 11670 11396 11726 11398
rect 11750 11396 11806 11398
rect 15212 11450 15268 11452
rect 15292 11450 15348 11452
rect 15372 11450 15428 11452
rect 15452 11450 15508 11452
rect 15212 11398 15258 11450
rect 15258 11398 15268 11450
rect 15292 11398 15322 11450
rect 15322 11398 15334 11450
rect 15334 11398 15348 11450
rect 15372 11398 15386 11450
rect 15386 11398 15398 11450
rect 15398 11398 15428 11450
rect 15452 11398 15462 11450
rect 15462 11398 15508 11450
rect 15212 11396 15268 11398
rect 15292 11396 15348 11398
rect 15372 11396 15428 11398
rect 15452 11396 15508 11398
rect 13361 10906 13417 10908
rect 13441 10906 13497 10908
rect 13521 10906 13577 10908
rect 13601 10906 13657 10908
rect 13361 10854 13407 10906
rect 13407 10854 13417 10906
rect 13441 10854 13471 10906
rect 13471 10854 13483 10906
rect 13483 10854 13497 10906
rect 13521 10854 13535 10906
rect 13535 10854 13547 10906
rect 13547 10854 13577 10906
rect 13601 10854 13611 10906
rect 13611 10854 13657 10906
rect 13361 10852 13417 10854
rect 13441 10852 13497 10854
rect 13521 10852 13577 10854
rect 13601 10852 13657 10854
rect 11510 10362 11566 10364
rect 11590 10362 11646 10364
rect 11670 10362 11726 10364
rect 11750 10362 11806 10364
rect 11510 10310 11556 10362
rect 11556 10310 11566 10362
rect 11590 10310 11620 10362
rect 11620 10310 11632 10362
rect 11632 10310 11646 10362
rect 11670 10310 11684 10362
rect 11684 10310 11696 10362
rect 11696 10310 11726 10362
rect 11750 10310 11760 10362
rect 11760 10310 11806 10362
rect 11510 10308 11566 10310
rect 11590 10308 11646 10310
rect 11670 10308 11726 10310
rect 11750 10308 11806 10310
rect 15212 10362 15268 10364
rect 15292 10362 15348 10364
rect 15372 10362 15428 10364
rect 15452 10362 15508 10364
rect 15212 10310 15258 10362
rect 15258 10310 15268 10362
rect 15292 10310 15322 10362
rect 15322 10310 15334 10362
rect 15334 10310 15348 10362
rect 15372 10310 15386 10362
rect 15386 10310 15398 10362
rect 15398 10310 15428 10362
rect 15452 10310 15462 10362
rect 15462 10310 15508 10362
rect 15212 10308 15268 10310
rect 15292 10308 15348 10310
rect 15372 10308 15428 10310
rect 15452 10308 15508 10310
rect 13361 9818 13417 9820
rect 13441 9818 13497 9820
rect 13521 9818 13577 9820
rect 13601 9818 13657 9820
rect 13361 9766 13407 9818
rect 13407 9766 13417 9818
rect 13441 9766 13471 9818
rect 13471 9766 13483 9818
rect 13483 9766 13497 9818
rect 13521 9766 13535 9818
rect 13535 9766 13547 9818
rect 13547 9766 13577 9818
rect 13601 9766 13611 9818
rect 13611 9766 13657 9818
rect 13361 9764 13417 9766
rect 13441 9764 13497 9766
rect 13521 9764 13577 9766
rect 13601 9764 13657 9766
rect 11510 9274 11566 9276
rect 11590 9274 11646 9276
rect 11670 9274 11726 9276
rect 11750 9274 11806 9276
rect 11510 9222 11556 9274
rect 11556 9222 11566 9274
rect 11590 9222 11620 9274
rect 11620 9222 11632 9274
rect 11632 9222 11646 9274
rect 11670 9222 11684 9274
rect 11684 9222 11696 9274
rect 11696 9222 11726 9274
rect 11750 9222 11760 9274
rect 11760 9222 11806 9274
rect 11510 9220 11566 9222
rect 11590 9220 11646 9222
rect 11670 9220 11726 9222
rect 11750 9220 11806 9222
rect 15212 9274 15268 9276
rect 15292 9274 15348 9276
rect 15372 9274 15428 9276
rect 15452 9274 15508 9276
rect 15212 9222 15258 9274
rect 15258 9222 15268 9274
rect 15292 9222 15322 9274
rect 15322 9222 15334 9274
rect 15334 9222 15348 9274
rect 15372 9222 15386 9274
rect 15386 9222 15398 9274
rect 15398 9222 15428 9274
rect 15452 9222 15462 9274
rect 15462 9222 15508 9274
rect 15212 9220 15268 9222
rect 15292 9220 15348 9222
rect 15372 9220 15428 9222
rect 15452 9220 15508 9222
rect 13361 8730 13417 8732
rect 13441 8730 13497 8732
rect 13521 8730 13577 8732
rect 13601 8730 13657 8732
rect 13361 8678 13407 8730
rect 13407 8678 13417 8730
rect 13441 8678 13471 8730
rect 13471 8678 13483 8730
rect 13483 8678 13497 8730
rect 13521 8678 13535 8730
rect 13535 8678 13547 8730
rect 13547 8678 13577 8730
rect 13601 8678 13611 8730
rect 13611 8678 13657 8730
rect 13361 8676 13417 8678
rect 13441 8676 13497 8678
rect 13521 8676 13577 8678
rect 13601 8676 13657 8678
rect 11510 8186 11566 8188
rect 11590 8186 11646 8188
rect 11670 8186 11726 8188
rect 11750 8186 11806 8188
rect 11510 8134 11556 8186
rect 11556 8134 11566 8186
rect 11590 8134 11620 8186
rect 11620 8134 11632 8186
rect 11632 8134 11646 8186
rect 11670 8134 11684 8186
rect 11684 8134 11696 8186
rect 11696 8134 11726 8186
rect 11750 8134 11760 8186
rect 11760 8134 11806 8186
rect 11510 8132 11566 8134
rect 11590 8132 11646 8134
rect 11670 8132 11726 8134
rect 11750 8132 11806 8134
rect 15212 8186 15268 8188
rect 15292 8186 15348 8188
rect 15372 8186 15428 8188
rect 15452 8186 15508 8188
rect 15212 8134 15258 8186
rect 15258 8134 15268 8186
rect 15292 8134 15322 8186
rect 15322 8134 15334 8186
rect 15334 8134 15348 8186
rect 15372 8134 15386 8186
rect 15386 8134 15398 8186
rect 15398 8134 15428 8186
rect 15452 8134 15462 8186
rect 15462 8134 15508 8186
rect 15212 8132 15268 8134
rect 15292 8132 15348 8134
rect 15372 8132 15428 8134
rect 15452 8132 15508 8134
rect 13361 7642 13417 7644
rect 13441 7642 13497 7644
rect 13521 7642 13577 7644
rect 13601 7642 13657 7644
rect 13361 7590 13407 7642
rect 13407 7590 13417 7642
rect 13441 7590 13471 7642
rect 13471 7590 13483 7642
rect 13483 7590 13497 7642
rect 13521 7590 13535 7642
rect 13535 7590 13547 7642
rect 13547 7590 13577 7642
rect 13601 7590 13611 7642
rect 13611 7590 13657 7642
rect 13361 7588 13417 7590
rect 13441 7588 13497 7590
rect 13521 7588 13577 7590
rect 13601 7588 13657 7590
rect 11510 7098 11566 7100
rect 11590 7098 11646 7100
rect 11670 7098 11726 7100
rect 11750 7098 11806 7100
rect 11510 7046 11556 7098
rect 11556 7046 11566 7098
rect 11590 7046 11620 7098
rect 11620 7046 11632 7098
rect 11632 7046 11646 7098
rect 11670 7046 11684 7098
rect 11684 7046 11696 7098
rect 11696 7046 11726 7098
rect 11750 7046 11760 7098
rect 11760 7046 11806 7098
rect 11510 7044 11566 7046
rect 11590 7044 11646 7046
rect 11670 7044 11726 7046
rect 11750 7044 11806 7046
rect 15212 7098 15268 7100
rect 15292 7098 15348 7100
rect 15372 7098 15428 7100
rect 15452 7098 15508 7100
rect 15212 7046 15258 7098
rect 15258 7046 15268 7098
rect 15292 7046 15322 7098
rect 15322 7046 15334 7098
rect 15334 7046 15348 7098
rect 15372 7046 15386 7098
rect 15386 7046 15398 7098
rect 15398 7046 15428 7098
rect 15452 7046 15462 7098
rect 15462 7046 15508 7098
rect 15212 7044 15268 7046
rect 15292 7044 15348 7046
rect 15372 7044 15428 7046
rect 15452 7044 15508 7046
rect 2255 6554 2311 6556
rect 2335 6554 2391 6556
rect 2415 6554 2471 6556
rect 2495 6554 2551 6556
rect 2255 6502 2301 6554
rect 2301 6502 2311 6554
rect 2335 6502 2365 6554
rect 2365 6502 2377 6554
rect 2377 6502 2391 6554
rect 2415 6502 2429 6554
rect 2429 6502 2441 6554
rect 2441 6502 2471 6554
rect 2495 6502 2505 6554
rect 2505 6502 2551 6554
rect 2255 6500 2311 6502
rect 2335 6500 2391 6502
rect 2415 6500 2471 6502
rect 2495 6500 2551 6502
rect 5957 6554 6013 6556
rect 6037 6554 6093 6556
rect 6117 6554 6173 6556
rect 6197 6554 6253 6556
rect 5957 6502 6003 6554
rect 6003 6502 6013 6554
rect 6037 6502 6067 6554
rect 6067 6502 6079 6554
rect 6079 6502 6093 6554
rect 6117 6502 6131 6554
rect 6131 6502 6143 6554
rect 6143 6502 6173 6554
rect 6197 6502 6207 6554
rect 6207 6502 6253 6554
rect 5957 6500 6013 6502
rect 6037 6500 6093 6502
rect 6117 6500 6173 6502
rect 6197 6500 6253 6502
rect 9659 6554 9715 6556
rect 9739 6554 9795 6556
rect 9819 6554 9875 6556
rect 9899 6554 9955 6556
rect 9659 6502 9705 6554
rect 9705 6502 9715 6554
rect 9739 6502 9769 6554
rect 9769 6502 9781 6554
rect 9781 6502 9795 6554
rect 9819 6502 9833 6554
rect 9833 6502 9845 6554
rect 9845 6502 9875 6554
rect 9899 6502 9909 6554
rect 9909 6502 9955 6554
rect 9659 6500 9715 6502
rect 9739 6500 9795 6502
rect 9819 6500 9875 6502
rect 9899 6500 9955 6502
rect 4106 6010 4162 6012
rect 4186 6010 4242 6012
rect 4266 6010 4322 6012
rect 4346 6010 4402 6012
rect 4106 5958 4152 6010
rect 4152 5958 4162 6010
rect 4186 5958 4216 6010
rect 4216 5958 4228 6010
rect 4228 5958 4242 6010
rect 4266 5958 4280 6010
rect 4280 5958 4292 6010
rect 4292 5958 4322 6010
rect 4346 5958 4356 6010
rect 4356 5958 4402 6010
rect 4106 5956 4162 5958
rect 4186 5956 4242 5958
rect 4266 5956 4322 5958
rect 4346 5956 4402 5958
rect 7808 6010 7864 6012
rect 7888 6010 7944 6012
rect 7968 6010 8024 6012
rect 8048 6010 8104 6012
rect 7808 5958 7854 6010
rect 7854 5958 7864 6010
rect 7888 5958 7918 6010
rect 7918 5958 7930 6010
rect 7930 5958 7944 6010
rect 7968 5958 7982 6010
rect 7982 5958 7994 6010
rect 7994 5958 8024 6010
rect 8048 5958 8058 6010
rect 8058 5958 8104 6010
rect 7808 5956 7864 5958
rect 7888 5956 7944 5958
rect 7968 5956 8024 5958
rect 8048 5956 8104 5958
rect 2255 5466 2311 5468
rect 2335 5466 2391 5468
rect 2415 5466 2471 5468
rect 2495 5466 2551 5468
rect 2255 5414 2301 5466
rect 2301 5414 2311 5466
rect 2335 5414 2365 5466
rect 2365 5414 2377 5466
rect 2377 5414 2391 5466
rect 2415 5414 2429 5466
rect 2429 5414 2441 5466
rect 2441 5414 2471 5466
rect 2495 5414 2505 5466
rect 2505 5414 2551 5466
rect 2255 5412 2311 5414
rect 2335 5412 2391 5414
rect 2415 5412 2471 5414
rect 2495 5412 2551 5414
rect 5957 5466 6013 5468
rect 6037 5466 6093 5468
rect 6117 5466 6173 5468
rect 6197 5466 6253 5468
rect 5957 5414 6003 5466
rect 6003 5414 6013 5466
rect 6037 5414 6067 5466
rect 6067 5414 6079 5466
rect 6079 5414 6093 5466
rect 6117 5414 6131 5466
rect 6131 5414 6143 5466
rect 6143 5414 6173 5466
rect 6197 5414 6207 5466
rect 6207 5414 6253 5466
rect 5957 5412 6013 5414
rect 6037 5412 6093 5414
rect 6117 5412 6173 5414
rect 6197 5412 6253 5414
rect 9659 5466 9715 5468
rect 9739 5466 9795 5468
rect 9819 5466 9875 5468
rect 9899 5466 9955 5468
rect 9659 5414 9705 5466
rect 9705 5414 9715 5466
rect 9739 5414 9769 5466
rect 9769 5414 9781 5466
rect 9781 5414 9795 5466
rect 9819 5414 9833 5466
rect 9833 5414 9845 5466
rect 9845 5414 9875 5466
rect 9899 5414 9909 5466
rect 9909 5414 9955 5466
rect 9659 5412 9715 5414
rect 9739 5412 9795 5414
rect 9819 5412 9875 5414
rect 9899 5412 9955 5414
rect 4106 4922 4162 4924
rect 4186 4922 4242 4924
rect 4266 4922 4322 4924
rect 4346 4922 4402 4924
rect 4106 4870 4152 4922
rect 4152 4870 4162 4922
rect 4186 4870 4216 4922
rect 4216 4870 4228 4922
rect 4228 4870 4242 4922
rect 4266 4870 4280 4922
rect 4280 4870 4292 4922
rect 4292 4870 4322 4922
rect 4346 4870 4356 4922
rect 4356 4870 4402 4922
rect 4106 4868 4162 4870
rect 4186 4868 4242 4870
rect 4266 4868 4322 4870
rect 4346 4868 4402 4870
rect 7808 4922 7864 4924
rect 7888 4922 7944 4924
rect 7968 4922 8024 4924
rect 8048 4922 8104 4924
rect 7808 4870 7854 4922
rect 7854 4870 7864 4922
rect 7888 4870 7918 4922
rect 7918 4870 7930 4922
rect 7930 4870 7944 4922
rect 7968 4870 7982 4922
rect 7982 4870 7994 4922
rect 7994 4870 8024 4922
rect 8048 4870 8058 4922
rect 8058 4870 8104 4922
rect 7808 4868 7864 4870
rect 7888 4868 7944 4870
rect 7968 4868 8024 4870
rect 8048 4868 8104 4870
rect 13361 6554 13417 6556
rect 13441 6554 13497 6556
rect 13521 6554 13577 6556
rect 13601 6554 13657 6556
rect 13361 6502 13407 6554
rect 13407 6502 13417 6554
rect 13441 6502 13471 6554
rect 13471 6502 13483 6554
rect 13483 6502 13497 6554
rect 13521 6502 13535 6554
rect 13535 6502 13547 6554
rect 13547 6502 13577 6554
rect 13601 6502 13611 6554
rect 13611 6502 13657 6554
rect 13361 6500 13417 6502
rect 13441 6500 13497 6502
rect 13521 6500 13577 6502
rect 13601 6500 13657 6502
rect 11510 6010 11566 6012
rect 11590 6010 11646 6012
rect 11670 6010 11726 6012
rect 11750 6010 11806 6012
rect 11510 5958 11556 6010
rect 11556 5958 11566 6010
rect 11590 5958 11620 6010
rect 11620 5958 11632 6010
rect 11632 5958 11646 6010
rect 11670 5958 11684 6010
rect 11684 5958 11696 6010
rect 11696 5958 11726 6010
rect 11750 5958 11760 6010
rect 11760 5958 11806 6010
rect 11510 5956 11566 5958
rect 11590 5956 11646 5958
rect 11670 5956 11726 5958
rect 11750 5956 11806 5958
rect 15212 6010 15268 6012
rect 15292 6010 15348 6012
rect 15372 6010 15428 6012
rect 15452 6010 15508 6012
rect 15212 5958 15258 6010
rect 15258 5958 15268 6010
rect 15292 5958 15322 6010
rect 15322 5958 15334 6010
rect 15334 5958 15348 6010
rect 15372 5958 15386 6010
rect 15386 5958 15398 6010
rect 15398 5958 15428 6010
rect 15452 5958 15462 6010
rect 15462 5958 15508 6010
rect 15212 5956 15268 5958
rect 15292 5956 15348 5958
rect 15372 5956 15428 5958
rect 15452 5956 15508 5958
rect 13361 5466 13417 5468
rect 13441 5466 13497 5468
rect 13521 5466 13577 5468
rect 13601 5466 13657 5468
rect 13361 5414 13407 5466
rect 13407 5414 13417 5466
rect 13441 5414 13471 5466
rect 13471 5414 13483 5466
rect 13483 5414 13497 5466
rect 13521 5414 13535 5466
rect 13535 5414 13547 5466
rect 13547 5414 13577 5466
rect 13601 5414 13611 5466
rect 13611 5414 13657 5466
rect 13361 5412 13417 5414
rect 13441 5412 13497 5414
rect 13521 5412 13577 5414
rect 13601 5412 13657 5414
rect 11510 4922 11566 4924
rect 11590 4922 11646 4924
rect 11670 4922 11726 4924
rect 11750 4922 11806 4924
rect 11510 4870 11556 4922
rect 11556 4870 11566 4922
rect 11590 4870 11620 4922
rect 11620 4870 11632 4922
rect 11632 4870 11646 4922
rect 11670 4870 11684 4922
rect 11684 4870 11696 4922
rect 11696 4870 11726 4922
rect 11750 4870 11760 4922
rect 11760 4870 11806 4922
rect 11510 4868 11566 4870
rect 11590 4868 11646 4870
rect 11670 4868 11726 4870
rect 11750 4868 11806 4870
rect 15212 4922 15268 4924
rect 15292 4922 15348 4924
rect 15372 4922 15428 4924
rect 15452 4922 15508 4924
rect 15212 4870 15258 4922
rect 15258 4870 15268 4922
rect 15292 4870 15322 4922
rect 15322 4870 15334 4922
rect 15334 4870 15348 4922
rect 15372 4870 15386 4922
rect 15386 4870 15398 4922
rect 15398 4870 15428 4922
rect 15452 4870 15462 4922
rect 15462 4870 15508 4922
rect 15212 4868 15268 4870
rect 15292 4868 15348 4870
rect 15372 4868 15428 4870
rect 15452 4868 15508 4870
rect 2255 4378 2311 4380
rect 2335 4378 2391 4380
rect 2415 4378 2471 4380
rect 2495 4378 2551 4380
rect 2255 4326 2301 4378
rect 2301 4326 2311 4378
rect 2335 4326 2365 4378
rect 2365 4326 2377 4378
rect 2377 4326 2391 4378
rect 2415 4326 2429 4378
rect 2429 4326 2441 4378
rect 2441 4326 2471 4378
rect 2495 4326 2505 4378
rect 2505 4326 2551 4378
rect 2255 4324 2311 4326
rect 2335 4324 2391 4326
rect 2415 4324 2471 4326
rect 2495 4324 2551 4326
rect 5957 4378 6013 4380
rect 6037 4378 6093 4380
rect 6117 4378 6173 4380
rect 6197 4378 6253 4380
rect 5957 4326 6003 4378
rect 6003 4326 6013 4378
rect 6037 4326 6067 4378
rect 6067 4326 6079 4378
rect 6079 4326 6093 4378
rect 6117 4326 6131 4378
rect 6131 4326 6143 4378
rect 6143 4326 6173 4378
rect 6197 4326 6207 4378
rect 6207 4326 6253 4378
rect 5957 4324 6013 4326
rect 6037 4324 6093 4326
rect 6117 4324 6173 4326
rect 6197 4324 6253 4326
rect 9659 4378 9715 4380
rect 9739 4378 9795 4380
rect 9819 4378 9875 4380
rect 9899 4378 9955 4380
rect 9659 4326 9705 4378
rect 9705 4326 9715 4378
rect 9739 4326 9769 4378
rect 9769 4326 9781 4378
rect 9781 4326 9795 4378
rect 9819 4326 9833 4378
rect 9833 4326 9845 4378
rect 9845 4326 9875 4378
rect 9899 4326 9909 4378
rect 9909 4326 9955 4378
rect 9659 4324 9715 4326
rect 9739 4324 9795 4326
rect 9819 4324 9875 4326
rect 9899 4324 9955 4326
rect 13361 4378 13417 4380
rect 13441 4378 13497 4380
rect 13521 4378 13577 4380
rect 13601 4378 13657 4380
rect 13361 4326 13407 4378
rect 13407 4326 13417 4378
rect 13441 4326 13471 4378
rect 13471 4326 13483 4378
rect 13483 4326 13497 4378
rect 13521 4326 13535 4378
rect 13535 4326 13547 4378
rect 13547 4326 13577 4378
rect 13601 4326 13611 4378
rect 13611 4326 13657 4378
rect 13361 4324 13417 4326
rect 13441 4324 13497 4326
rect 13521 4324 13577 4326
rect 13601 4324 13657 4326
rect 11242 4120 11298 4176
rect 4106 3834 4162 3836
rect 4186 3834 4242 3836
rect 4266 3834 4322 3836
rect 4346 3834 4402 3836
rect 4106 3782 4152 3834
rect 4152 3782 4162 3834
rect 4186 3782 4216 3834
rect 4216 3782 4228 3834
rect 4228 3782 4242 3834
rect 4266 3782 4280 3834
rect 4280 3782 4292 3834
rect 4292 3782 4322 3834
rect 4346 3782 4356 3834
rect 4356 3782 4402 3834
rect 4106 3780 4162 3782
rect 4186 3780 4242 3782
rect 4266 3780 4322 3782
rect 4346 3780 4402 3782
rect 7808 3834 7864 3836
rect 7888 3834 7944 3836
rect 7968 3834 8024 3836
rect 8048 3834 8104 3836
rect 7808 3782 7854 3834
rect 7854 3782 7864 3834
rect 7888 3782 7918 3834
rect 7918 3782 7930 3834
rect 7930 3782 7944 3834
rect 7968 3782 7982 3834
rect 7982 3782 7994 3834
rect 7994 3782 8024 3834
rect 8048 3782 8058 3834
rect 8058 3782 8104 3834
rect 7808 3780 7864 3782
rect 7888 3780 7944 3782
rect 7968 3780 8024 3782
rect 8048 3780 8104 3782
rect 11510 3834 11566 3836
rect 11590 3834 11646 3836
rect 11670 3834 11726 3836
rect 11750 3834 11806 3836
rect 11510 3782 11556 3834
rect 11556 3782 11566 3834
rect 11590 3782 11620 3834
rect 11620 3782 11632 3834
rect 11632 3782 11646 3834
rect 11670 3782 11684 3834
rect 11684 3782 11696 3834
rect 11696 3782 11726 3834
rect 11750 3782 11760 3834
rect 11760 3782 11806 3834
rect 11510 3780 11566 3782
rect 11590 3780 11646 3782
rect 11670 3780 11726 3782
rect 11750 3780 11806 3782
rect 15212 3834 15268 3836
rect 15292 3834 15348 3836
rect 15372 3834 15428 3836
rect 15452 3834 15508 3836
rect 15212 3782 15258 3834
rect 15258 3782 15268 3834
rect 15292 3782 15322 3834
rect 15322 3782 15334 3834
rect 15334 3782 15348 3834
rect 15372 3782 15386 3834
rect 15386 3782 15398 3834
rect 15398 3782 15428 3834
rect 15452 3782 15462 3834
rect 15462 3782 15508 3834
rect 15212 3780 15268 3782
rect 15292 3780 15348 3782
rect 15372 3780 15428 3782
rect 15452 3780 15508 3782
rect 2255 3290 2311 3292
rect 2335 3290 2391 3292
rect 2415 3290 2471 3292
rect 2495 3290 2551 3292
rect 2255 3238 2301 3290
rect 2301 3238 2311 3290
rect 2335 3238 2365 3290
rect 2365 3238 2377 3290
rect 2377 3238 2391 3290
rect 2415 3238 2429 3290
rect 2429 3238 2441 3290
rect 2441 3238 2471 3290
rect 2495 3238 2505 3290
rect 2505 3238 2551 3290
rect 2255 3236 2311 3238
rect 2335 3236 2391 3238
rect 2415 3236 2471 3238
rect 2495 3236 2551 3238
rect 5957 3290 6013 3292
rect 6037 3290 6093 3292
rect 6117 3290 6173 3292
rect 6197 3290 6253 3292
rect 5957 3238 6003 3290
rect 6003 3238 6013 3290
rect 6037 3238 6067 3290
rect 6067 3238 6079 3290
rect 6079 3238 6093 3290
rect 6117 3238 6131 3290
rect 6131 3238 6143 3290
rect 6143 3238 6173 3290
rect 6197 3238 6207 3290
rect 6207 3238 6253 3290
rect 5957 3236 6013 3238
rect 6037 3236 6093 3238
rect 6117 3236 6173 3238
rect 6197 3236 6253 3238
rect 9659 3290 9715 3292
rect 9739 3290 9795 3292
rect 9819 3290 9875 3292
rect 9899 3290 9955 3292
rect 9659 3238 9705 3290
rect 9705 3238 9715 3290
rect 9739 3238 9769 3290
rect 9769 3238 9781 3290
rect 9781 3238 9795 3290
rect 9819 3238 9833 3290
rect 9833 3238 9845 3290
rect 9845 3238 9875 3290
rect 9899 3238 9909 3290
rect 9909 3238 9955 3290
rect 9659 3236 9715 3238
rect 9739 3236 9795 3238
rect 9819 3236 9875 3238
rect 9899 3236 9955 3238
rect 13361 3290 13417 3292
rect 13441 3290 13497 3292
rect 13521 3290 13577 3292
rect 13601 3290 13657 3292
rect 13361 3238 13407 3290
rect 13407 3238 13417 3290
rect 13441 3238 13471 3290
rect 13471 3238 13483 3290
rect 13483 3238 13497 3290
rect 13521 3238 13535 3290
rect 13535 3238 13547 3290
rect 13547 3238 13577 3290
rect 13601 3238 13611 3290
rect 13611 3238 13657 3290
rect 13361 3236 13417 3238
rect 13441 3236 13497 3238
rect 13521 3236 13577 3238
rect 13601 3236 13657 3238
rect 4106 2746 4162 2748
rect 4186 2746 4242 2748
rect 4266 2746 4322 2748
rect 4346 2746 4402 2748
rect 4106 2694 4152 2746
rect 4152 2694 4162 2746
rect 4186 2694 4216 2746
rect 4216 2694 4228 2746
rect 4228 2694 4242 2746
rect 4266 2694 4280 2746
rect 4280 2694 4292 2746
rect 4292 2694 4322 2746
rect 4346 2694 4356 2746
rect 4356 2694 4402 2746
rect 4106 2692 4162 2694
rect 4186 2692 4242 2694
rect 4266 2692 4322 2694
rect 4346 2692 4402 2694
rect 7808 2746 7864 2748
rect 7888 2746 7944 2748
rect 7968 2746 8024 2748
rect 8048 2746 8104 2748
rect 7808 2694 7854 2746
rect 7854 2694 7864 2746
rect 7888 2694 7918 2746
rect 7918 2694 7930 2746
rect 7930 2694 7944 2746
rect 7968 2694 7982 2746
rect 7982 2694 7994 2746
rect 7994 2694 8024 2746
rect 8048 2694 8058 2746
rect 8058 2694 8104 2746
rect 7808 2692 7864 2694
rect 7888 2692 7944 2694
rect 7968 2692 8024 2694
rect 8048 2692 8104 2694
rect 11510 2746 11566 2748
rect 11590 2746 11646 2748
rect 11670 2746 11726 2748
rect 11750 2746 11806 2748
rect 11510 2694 11556 2746
rect 11556 2694 11566 2746
rect 11590 2694 11620 2746
rect 11620 2694 11632 2746
rect 11632 2694 11646 2746
rect 11670 2694 11684 2746
rect 11684 2694 11696 2746
rect 11696 2694 11726 2746
rect 11750 2694 11760 2746
rect 11760 2694 11806 2746
rect 11510 2692 11566 2694
rect 11590 2692 11646 2694
rect 11670 2692 11726 2694
rect 11750 2692 11806 2694
rect 15212 2746 15268 2748
rect 15292 2746 15348 2748
rect 15372 2746 15428 2748
rect 15452 2746 15508 2748
rect 15212 2694 15258 2746
rect 15258 2694 15268 2746
rect 15292 2694 15322 2746
rect 15322 2694 15334 2746
rect 15334 2694 15348 2746
rect 15372 2694 15386 2746
rect 15386 2694 15398 2746
rect 15398 2694 15428 2746
rect 15452 2694 15462 2746
rect 15462 2694 15508 2746
rect 15212 2692 15268 2694
rect 15292 2692 15348 2694
rect 15372 2692 15428 2694
rect 15452 2692 15508 2694
rect 2255 2202 2311 2204
rect 2335 2202 2391 2204
rect 2415 2202 2471 2204
rect 2495 2202 2551 2204
rect 2255 2150 2301 2202
rect 2301 2150 2311 2202
rect 2335 2150 2365 2202
rect 2365 2150 2377 2202
rect 2377 2150 2391 2202
rect 2415 2150 2429 2202
rect 2429 2150 2441 2202
rect 2441 2150 2471 2202
rect 2495 2150 2505 2202
rect 2505 2150 2551 2202
rect 2255 2148 2311 2150
rect 2335 2148 2391 2150
rect 2415 2148 2471 2150
rect 2495 2148 2551 2150
rect 5957 2202 6013 2204
rect 6037 2202 6093 2204
rect 6117 2202 6173 2204
rect 6197 2202 6253 2204
rect 5957 2150 6003 2202
rect 6003 2150 6013 2202
rect 6037 2150 6067 2202
rect 6067 2150 6079 2202
rect 6079 2150 6093 2202
rect 6117 2150 6131 2202
rect 6131 2150 6143 2202
rect 6143 2150 6173 2202
rect 6197 2150 6207 2202
rect 6207 2150 6253 2202
rect 5957 2148 6013 2150
rect 6037 2148 6093 2150
rect 6117 2148 6173 2150
rect 6197 2148 6253 2150
rect 9659 2202 9715 2204
rect 9739 2202 9795 2204
rect 9819 2202 9875 2204
rect 9899 2202 9955 2204
rect 9659 2150 9705 2202
rect 9705 2150 9715 2202
rect 9739 2150 9769 2202
rect 9769 2150 9781 2202
rect 9781 2150 9795 2202
rect 9819 2150 9833 2202
rect 9833 2150 9845 2202
rect 9845 2150 9875 2202
rect 9899 2150 9909 2202
rect 9909 2150 9955 2202
rect 9659 2148 9715 2150
rect 9739 2148 9795 2150
rect 9819 2148 9875 2150
rect 9899 2148 9955 2150
rect 13361 2202 13417 2204
rect 13441 2202 13497 2204
rect 13521 2202 13577 2204
rect 13601 2202 13657 2204
rect 13361 2150 13407 2202
rect 13407 2150 13417 2202
rect 13441 2150 13471 2202
rect 13471 2150 13483 2202
rect 13483 2150 13497 2202
rect 13521 2150 13535 2202
rect 13535 2150 13547 2202
rect 13547 2150 13577 2202
rect 13601 2150 13611 2202
rect 13611 2150 13657 2202
rect 13361 2148 13417 2150
rect 13441 2148 13497 2150
rect 13521 2148 13577 2150
rect 13601 2148 13657 2150
rect 4106 1658 4162 1660
rect 4186 1658 4242 1660
rect 4266 1658 4322 1660
rect 4346 1658 4402 1660
rect 4106 1606 4152 1658
rect 4152 1606 4162 1658
rect 4186 1606 4216 1658
rect 4216 1606 4228 1658
rect 4228 1606 4242 1658
rect 4266 1606 4280 1658
rect 4280 1606 4292 1658
rect 4292 1606 4322 1658
rect 4346 1606 4356 1658
rect 4356 1606 4402 1658
rect 4106 1604 4162 1606
rect 4186 1604 4242 1606
rect 4266 1604 4322 1606
rect 4346 1604 4402 1606
rect 7808 1658 7864 1660
rect 7888 1658 7944 1660
rect 7968 1658 8024 1660
rect 8048 1658 8104 1660
rect 7808 1606 7854 1658
rect 7854 1606 7864 1658
rect 7888 1606 7918 1658
rect 7918 1606 7930 1658
rect 7930 1606 7944 1658
rect 7968 1606 7982 1658
rect 7982 1606 7994 1658
rect 7994 1606 8024 1658
rect 8048 1606 8058 1658
rect 8058 1606 8104 1658
rect 7808 1604 7864 1606
rect 7888 1604 7944 1606
rect 7968 1604 8024 1606
rect 8048 1604 8104 1606
rect 11510 1658 11566 1660
rect 11590 1658 11646 1660
rect 11670 1658 11726 1660
rect 11750 1658 11806 1660
rect 11510 1606 11556 1658
rect 11556 1606 11566 1658
rect 11590 1606 11620 1658
rect 11620 1606 11632 1658
rect 11632 1606 11646 1658
rect 11670 1606 11684 1658
rect 11684 1606 11696 1658
rect 11696 1606 11726 1658
rect 11750 1606 11760 1658
rect 11760 1606 11806 1658
rect 11510 1604 11566 1606
rect 11590 1604 11646 1606
rect 11670 1604 11726 1606
rect 11750 1604 11806 1606
rect 15212 1658 15268 1660
rect 15292 1658 15348 1660
rect 15372 1658 15428 1660
rect 15452 1658 15508 1660
rect 15212 1606 15258 1658
rect 15258 1606 15268 1658
rect 15292 1606 15322 1658
rect 15322 1606 15334 1658
rect 15334 1606 15348 1658
rect 15372 1606 15386 1658
rect 15386 1606 15398 1658
rect 15398 1606 15428 1658
rect 15452 1606 15462 1658
rect 15462 1606 15508 1658
rect 15212 1604 15268 1606
rect 15292 1604 15348 1606
rect 15372 1604 15428 1606
rect 15452 1604 15508 1606
rect 2255 1114 2311 1116
rect 2335 1114 2391 1116
rect 2415 1114 2471 1116
rect 2495 1114 2551 1116
rect 2255 1062 2301 1114
rect 2301 1062 2311 1114
rect 2335 1062 2365 1114
rect 2365 1062 2377 1114
rect 2377 1062 2391 1114
rect 2415 1062 2429 1114
rect 2429 1062 2441 1114
rect 2441 1062 2471 1114
rect 2495 1062 2505 1114
rect 2505 1062 2551 1114
rect 2255 1060 2311 1062
rect 2335 1060 2391 1062
rect 2415 1060 2471 1062
rect 2495 1060 2551 1062
rect 5957 1114 6013 1116
rect 6037 1114 6093 1116
rect 6117 1114 6173 1116
rect 6197 1114 6253 1116
rect 5957 1062 6003 1114
rect 6003 1062 6013 1114
rect 6037 1062 6067 1114
rect 6067 1062 6079 1114
rect 6079 1062 6093 1114
rect 6117 1062 6131 1114
rect 6131 1062 6143 1114
rect 6143 1062 6173 1114
rect 6197 1062 6207 1114
rect 6207 1062 6253 1114
rect 5957 1060 6013 1062
rect 6037 1060 6093 1062
rect 6117 1060 6173 1062
rect 6197 1060 6253 1062
rect 9659 1114 9715 1116
rect 9739 1114 9795 1116
rect 9819 1114 9875 1116
rect 9899 1114 9955 1116
rect 9659 1062 9705 1114
rect 9705 1062 9715 1114
rect 9739 1062 9769 1114
rect 9769 1062 9781 1114
rect 9781 1062 9795 1114
rect 9819 1062 9833 1114
rect 9833 1062 9845 1114
rect 9845 1062 9875 1114
rect 9899 1062 9909 1114
rect 9909 1062 9955 1114
rect 9659 1060 9715 1062
rect 9739 1060 9795 1062
rect 9819 1060 9875 1062
rect 9899 1060 9955 1062
rect 13361 1114 13417 1116
rect 13441 1114 13497 1116
rect 13521 1114 13577 1116
rect 13601 1114 13657 1116
rect 13361 1062 13407 1114
rect 13407 1062 13417 1114
rect 13441 1062 13471 1114
rect 13471 1062 13483 1114
rect 13483 1062 13497 1114
rect 13521 1062 13535 1114
rect 13535 1062 13547 1114
rect 13547 1062 13577 1114
rect 13601 1062 13611 1114
rect 13611 1062 13657 1114
rect 13361 1060 13417 1062
rect 13441 1060 13497 1062
rect 13521 1060 13577 1062
rect 13601 1060 13657 1062
rect 4106 570 4162 572
rect 4186 570 4242 572
rect 4266 570 4322 572
rect 4346 570 4402 572
rect 4106 518 4152 570
rect 4152 518 4162 570
rect 4186 518 4216 570
rect 4216 518 4228 570
rect 4228 518 4242 570
rect 4266 518 4280 570
rect 4280 518 4292 570
rect 4292 518 4322 570
rect 4346 518 4356 570
rect 4356 518 4402 570
rect 4106 516 4162 518
rect 4186 516 4242 518
rect 4266 516 4322 518
rect 4346 516 4402 518
rect 7808 570 7864 572
rect 7888 570 7944 572
rect 7968 570 8024 572
rect 8048 570 8104 572
rect 7808 518 7854 570
rect 7854 518 7864 570
rect 7888 518 7918 570
rect 7918 518 7930 570
rect 7930 518 7944 570
rect 7968 518 7982 570
rect 7982 518 7994 570
rect 7994 518 8024 570
rect 8048 518 8058 570
rect 8058 518 8104 570
rect 7808 516 7864 518
rect 7888 516 7944 518
rect 7968 516 8024 518
rect 8048 516 8104 518
rect 11510 570 11566 572
rect 11590 570 11646 572
rect 11670 570 11726 572
rect 11750 570 11806 572
rect 11510 518 11556 570
rect 11556 518 11566 570
rect 11590 518 11620 570
rect 11620 518 11632 570
rect 11632 518 11646 570
rect 11670 518 11684 570
rect 11684 518 11696 570
rect 11696 518 11726 570
rect 11750 518 11760 570
rect 11760 518 11806 570
rect 11510 516 11566 518
rect 11590 516 11646 518
rect 11670 516 11726 518
rect 11750 516 11806 518
rect 15212 570 15268 572
rect 15292 570 15348 572
rect 15372 570 15428 572
rect 15452 570 15508 572
rect 15212 518 15258 570
rect 15258 518 15268 570
rect 15292 518 15322 570
rect 15322 518 15334 570
rect 15334 518 15348 570
rect 15372 518 15386 570
rect 15386 518 15398 570
rect 15398 518 15428 570
rect 15452 518 15462 570
rect 15462 518 15508 570
rect 15212 516 15268 518
rect 15292 516 15348 518
rect 15372 516 15428 518
rect 15452 516 15508 518
<< metal3 >>
rect 2245 15264 2561 15265
rect 2245 15200 2251 15264
rect 2315 15200 2331 15264
rect 2395 15200 2411 15264
rect 2475 15200 2491 15264
rect 2555 15200 2561 15264
rect 2245 15199 2561 15200
rect 5947 15264 6263 15265
rect 5947 15200 5953 15264
rect 6017 15200 6033 15264
rect 6097 15200 6113 15264
rect 6177 15200 6193 15264
rect 6257 15200 6263 15264
rect 5947 15199 6263 15200
rect 9649 15264 9965 15265
rect 9649 15200 9655 15264
rect 9719 15200 9735 15264
rect 9799 15200 9815 15264
rect 9879 15200 9895 15264
rect 9959 15200 9965 15264
rect 9649 15199 9965 15200
rect 13351 15264 13667 15265
rect 13351 15200 13357 15264
rect 13421 15200 13437 15264
rect 13501 15200 13517 15264
rect 13581 15200 13597 15264
rect 13661 15200 13667 15264
rect 13351 15199 13667 15200
rect 4096 14720 4412 14721
rect 4096 14656 4102 14720
rect 4166 14656 4182 14720
rect 4246 14656 4262 14720
rect 4326 14656 4342 14720
rect 4406 14656 4412 14720
rect 4096 14655 4412 14656
rect 7798 14720 8114 14721
rect 7798 14656 7804 14720
rect 7868 14656 7884 14720
rect 7948 14656 7964 14720
rect 8028 14656 8044 14720
rect 8108 14656 8114 14720
rect 7798 14655 8114 14656
rect 11500 14720 11816 14721
rect 11500 14656 11506 14720
rect 11570 14656 11586 14720
rect 11650 14656 11666 14720
rect 11730 14656 11746 14720
rect 11810 14656 11816 14720
rect 11500 14655 11816 14656
rect 15202 14720 15518 14721
rect 15202 14656 15208 14720
rect 15272 14656 15288 14720
rect 15352 14656 15368 14720
rect 15432 14656 15448 14720
rect 15512 14656 15518 14720
rect 15202 14655 15518 14656
rect 2245 14176 2561 14177
rect 2245 14112 2251 14176
rect 2315 14112 2331 14176
rect 2395 14112 2411 14176
rect 2475 14112 2491 14176
rect 2555 14112 2561 14176
rect 2245 14111 2561 14112
rect 5947 14176 6263 14177
rect 5947 14112 5953 14176
rect 6017 14112 6033 14176
rect 6097 14112 6113 14176
rect 6177 14112 6193 14176
rect 6257 14112 6263 14176
rect 5947 14111 6263 14112
rect 9649 14176 9965 14177
rect 9649 14112 9655 14176
rect 9719 14112 9735 14176
rect 9799 14112 9815 14176
rect 9879 14112 9895 14176
rect 9959 14112 9965 14176
rect 9649 14111 9965 14112
rect 13351 14176 13667 14177
rect 13351 14112 13357 14176
rect 13421 14112 13437 14176
rect 13501 14112 13517 14176
rect 13581 14112 13597 14176
rect 13661 14112 13667 14176
rect 13351 14111 13667 14112
rect 4096 13632 4412 13633
rect 4096 13568 4102 13632
rect 4166 13568 4182 13632
rect 4246 13568 4262 13632
rect 4326 13568 4342 13632
rect 4406 13568 4412 13632
rect 4096 13567 4412 13568
rect 7798 13632 8114 13633
rect 7798 13568 7804 13632
rect 7868 13568 7884 13632
rect 7948 13568 7964 13632
rect 8028 13568 8044 13632
rect 8108 13568 8114 13632
rect 7798 13567 8114 13568
rect 11500 13632 11816 13633
rect 11500 13568 11506 13632
rect 11570 13568 11586 13632
rect 11650 13568 11666 13632
rect 11730 13568 11746 13632
rect 11810 13568 11816 13632
rect 11500 13567 11816 13568
rect 15202 13632 15518 13633
rect 15202 13568 15208 13632
rect 15272 13568 15288 13632
rect 15352 13568 15368 13632
rect 15432 13568 15448 13632
rect 15512 13568 15518 13632
rect 15202 13567 15518 13568
rect 2245 13088 2561 13089
rect 2245 13024 2251 13088
rect 2315 13024 2331 13088
rect 2395 13024 2411 13088
rect 2475 13024 2491 13088
rect 2555 13024 2561 13088
rect 2245 13023 2561 13024
rect 5947 13088 6263 13089
rect 5947 13024 5953 13088
rect 6017 13024 6033 13088
rect 6097 13024 6113 13088
rect 6177 13024 6193 13088
rect 6257 13024 6263 13088
rect 5947 13023 6263 13024
rect 9649 13088 9965 13089
rect 9649 13024 9655 13088
rect 9719 13024 9735 13088
rect 9799 13024 9815 13088
rect 9879 13024 9895 13088
rect 9959 13024 9965 13088
rect 9649 13023 9965 13024
rect 13351 13088 13667 13089
rect 13351 13024 13357 13088
rect 13421 13024 13437 13088
rect 13501 13024 13517 13088
rect 13581 13024 13597 13088
rect 13661 13024 13667 13088
rect 13351 13023 13667 13024
rect 4096 12544 4412 12545
rect 4096 12480 4102 12544
rect 4166 12480 4182 12544
rect 4246 12480 4262 12544
rect 4326 12480 4342 12544
rect 4406 12480 4412 12544
rect 4096 12479 4412 12480
rect 7798 12544 8114 12545
rect 7798 12480 7804 12544
rect 7868 12480 7884 12544
rect 7948 12480 7964 12544
rect 8028 12480 8044 12544
rect 8108 12480 8114 12544
rect 7798 12479 8114 12480
rect 11500 12544 11816 12545
rect 11500 12480 11506 12544
rect 11570 12480 11586 12544
rect 11650 12480 11666 12544
rect 11730 12480 11746 12544
rect 11810 12480 11816 12544
rect 11500 12479 11816 12480
rect 15202 12544 15518 12545
rect 15202 12480 15208 12544
rect 15272 12480 15288 12544
rect 15352 12480 15368 12544
rect 15432 12480 15448 12544
rect 15512 12480 15518 12544
rect 15202 12479 15518 12480
rect 2245 12000 2561 12001
rect 2245 11936 2251 12000
rect 2315 11936 2331 12000
rect 2395 11936 2411 12000
rect 2475 11936 2491 12000
rect 2555 11936 2561 12000
rect 2245 11935 2561 11936
rect 5947 12000 6263 12001
rect 5947 11936 5953 12000
rect 6017 11936 6033 12000
rect 6097 11936 6113 12000
rect 6177 11936 6193 12000
rect 6257 11936 6263 12000
rect 5947 11935 6263 11936
rect 9649 12000 9965 12001
rect 9649 11936 9655 12000
rect 9719 11936 9735 12000
rect 9799 11936 9815 12000
rect 9879 11936 9895 12000
rect 9959 11936 9965 12000
rect 9649 11935 9965 11936
rect 13351 12000 13667 12001
rect 13351 11936 13357 12000
rect 13421 11936 13437 12000
rect 13501 11936 13517 12000
rect 13581 11936 13597 12000
rect 13661 11936 13667 12000
rect 13351 11935 13667 11936
rect 14733 11794 14799 11797
rect 15600 11794 16000 11824
rect 14733 11792 16000 11794
rect 14733 11736 14738 11792
rect 14794 11736 16000 11792
rect 14733 11734 16000 11736
rect 14733 11731 14799 11734
rect 15600 11704 16000 11734
rect 4096 11456 4412 11457
rect 4096 11392 4102 11456
rect 4166 11392 4182 11456
rect 4246 11392 4262 11456
rect 4326 11392 4342 11456
rect 4406 11392 4412 11456
rect 4096 11391 4412 11392
rect 7798 11456 8114 11457
rect 7798 11392 7804 11456
rect 7868 11392 7884 11456
rect 7948 11392 7964 11456
rect 8028 11392 8044 11456
rect 8108 11392 8114 11456
rect 7798 11391 8114 11392
rect 11500 11456 11816 11457
rect 11500 11392 11506 11456
rect 11570 11392 11586 11456
rect 11650 11392 11666 11456
rect 11730 11392 11746 11456
rect 11810 11392 11816 11456
rect 11500 11391 11816 11392
rect 15202 11456 15518 11457
rect 15202 11392 15208 11456
rect 15272 11392 15288 11456
rect 15352 11392 15368 11456
rect 15432 11392 15448 11456
rect 15512 11392 15518 11456
rect 15202 11391 15518 11392
rect 2245 10912 2561 10913
rect 2245 10848 2251 10912
rect 2315 10848 2331 10912
rect 2395 10848 2411 10912
rect 2475 10848 2491 10912
rect 2555 10848 2561 10912
rect 2245 10847 2561 10848
rect 5947 10912 6263 10913
rect 5947 10848 5953 10912
rect 6017 10848 6033 10912
rect 6097 10848 6113 10912
rect 6177 10848 6193 10912
rect 6257 10848 6263 10912
rect 5947 10847 6263 10848
rect 9649 10912 9965 10913
rect 9649 10848 9655 10912
rect 9719 10848 9735 10912
rect 9799 10848 9815 10912
rect 9879 10848 9895 10912
rect 9959 10848 9965 10912
rect 9649 10847 9965 10848
rect 13351 10912 13667 10913
rect 13351 10848 13357 10912
rect 13421 10848 13437 10912
rect 13501 10848 13517 10912
rect 13581 10848 13597 10912
rect 13661 10848 13667 10912
rect 13351 10847 13667 10848
rect 4096 10368 4412 10369
rect 4096 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4342 10368
rect 4406 10304 4412 10368
rect 4096 10303 4412 10304
rect 7798 10368 8114 10369
rect 7798 10304 7804 10368
rect 7868 10304 7884 10368
rect 7948 10304 7964 10368
rect 8028 10304 8044 10368
rect 8108 10304 8114 10368
rect 7798 10303 8114 10304
rect 11500 10368 11816 10369
rect 11500 10304 11506 10368
rect 11570 10304 11586 10368
rect 11650 10304 11666 10368
rect 11730 10304 11746 10368
rect 11810 10304 11816 10368
rect 11500 10303 11816 10304
rect 15202 10368 15518 10369
rect 15202 10304 15208 10368
rect 15272 10304 15288 10368
rect 15352 10304 15368 10368
rect 15432 10304 15448 10368
rect 15512 10304 15518 10368
rect 15202 10303 15518 10304
rect 2245 9824 2561 9825
rect 2245 9760 2251 9824
rect 2315 9760 2331 9824
rect 2395 9760 2411 9824
rect 2475 9760 2491 9824
rect 2555 9760 2561 9824
rect 2245 9759 2561 9760
rect 5947 9824 6263 9825
rect 5947 9760 5953 9824
rect 6017 9760 6033 9824
rect 6097 9760 6113 9824
rect 6177 9760 6193 9824
rect 6257 9760 6263 9824
rect 5947 9759 6263 9760
rect 9649 9824 9965 9825
rect 9649 9760 9655 9824
rect 9719 9760 9735 9824
rect 9799 9760 9815 9824
rect 9879 9760 9895 9824
rect 9959 9760 9965 9824
rect 9649 9759 9965 9760
rect 13351 9824 13667 9825
rect 13351 9760 13357 9824
rect 13421 9760 13437 9824
rect 13501 9760 13517 9824
rect 13581 9760 13597 9824
rect 13661 9760 13667 9824
rect 13351 9759 13667 9760
rect 4096 9280 4412 9281
rect 4096 9216 4102 9280
rect 4166 9216 4182 9280
rect 4246 9216 4262 9280
rect 4326 9216 4342 9280
rect 4406 9216 4412 9280
rect 4096 9215 4412 9216
rect 7798 9280 8114 9281
rect 7798 9216 7804 9280
rect 7868 9216 7884 9280
rect 7948 9216 7964 9280
rect 8028 9216 8044 9280
rect 8108 9216 8114 9280
rect 7798 9215 8114 9216
rect 11500 9280 11816 9281
rect 11500 9216 11506 9280
rect 11570 9216 11586 9280
rect 11650 9216 11666 9280
rect 11730 9216 11746 9280
rect 11810 9216 11816 9280
rect 11500 9215 11816 9216
rect 15202 9280 15518 9281
rect 15202 9216 15208 9280
rect 15272 9216 15288 9280
rect 15352 9216 15368 9280
rect 15432 9216 15448 9280
rect 15512 9216 15518 9280
rect 15202 9215 15518 9216
rect 2245 8736 2561 8737
rect 2245 8672 2251 8736
rect 2315 8672 2331 8736
rect 2395 8672 2411 8736
rect 2475 8672 2491 8736
rect 2555 8672 2561 8736
rect 2245 8671 2561 8672
rect 5947 8736 6263 8737
rect 5947 8672 5953 8736
rect 6017 8672 6033 8736
rect 6097 8672 6113 8736
rect 6177 8672 6193 8736
rect 6257 8672 6263 8736
rect 5947 8671 6263 8672
rect 9649 8736 9965 8737
rect 9649 8672 9655 8736
rect 9719 8672 9735 8736
rect 9799 8672 9815 8736
rect 9879 8672 9895 8736
rect 9959 8672 9965 8736
rect 9649 8671 9965 8672
rect 13351 8736 13667 8737
rect 13351 8672 13357 8736
rect 13421 8672 13437 8736
rect 13501 8672 13517 8736
rect 13581 8672 13597 8736
rect 13661 8672 13667 8736
rect 13351 8671 13667 8672
rect 4096 8192 4412 8193
rect 4096 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4342 8192
rect 4406 8128 4412 8192
rect 4096 8127 4412 8128
rect 7798 8192 8114 8193
rect 7798 8128 7804 8192
rect 7868 8128 7884 8192
rect 7948 8128 7964 8192
rect 8028 8128 8044 8192
rect 8108 8128 8114 8192
rect 7798 8127 8114 8128
rect 11500 8192 11816 8193
rect 11500 8128 11506 8192
rect 11570 8128 11586 8192
rect 11650 8128 11666 8192
rect 11730 8128 11746 8192
rect 11810 8128 11816 8192
rect 11500 8127 11816 8128
rect 15202 8192 15518 8193
rect 15202 8128 15208 8192
rect 15272 8128 15288 8192
rect 15352 8128 15368 8192
rect 15432 8128 15448 8192
rect 15512 8128 15518 8192
rect 15202 8127 15518 8128
rect 2245 7648 2561 7649
rect 2245 7584 2251 7648
rect 2315 7584 2331 7648
rect 2395 7584 2411 7648
rect 2475 7584 2491 7648
rect 2555 7584 2561 7648
rect 2245 7583 2561 7584
rect 5947 7648 6263 7649
rect 5947 7584 5953 7648
rect 6017 7584 6033 7648
rect 6097 7584 6113 7648
rect 6177 7584 6193 7648
rect 6257 7584 6263 7648
rect 5947 7583 6263 7584
rect 9649 7648 9965 7649
rect 9649 7584 9655 7648
rect 9719 7584 9735 7648
rect 9799 7584 9815 7648
rect 9879 7584 9895 7648
rect 9959 7584 9965 7648
rect 9649 7583 9965 7584
rect 13351 7648 13667 7649
rect 13351 7584 13357 7648
rect 13421 7584 13437 7648
rect 13501 7584 13517 7648
rect 13581 7584 13597 7648
rect 13661 7584 13667 7648
rect 13351 7583 13667 7584
rect 4096 7104 4412 7105
rect 4096 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4342 7104
rect 4406 7040 4412 7104
rect 4096 7039 4412 7040
rect 7798 7104 8114 7105
rect 7798 7040 7804 7104
rect 7868 7040 7884 7104
rect 7948 7040 7964 7104
rect 8028 7040 8044 7104
rect 8108 7040 8114 7104
rect 7798 7039 8114 7040
rect 11500 7104 11816 7105
rect 11500 7040 11506 7104
rect 11570 7040 11586 7104
rect 11650 7040 11666 7104
rect 11730 7040 11746 7104
rect 11810 7040 11816 7104
rect 11500 7039 11816 7040
rect 15202 7104 15518 7105
rect 15202 7040 15208 7104
rect 15272 7040 15288 7104
rect 15352 7040 15368 7104
rect 15432 7040 15448 7104
rect 15512 7040 15518 7104
rect 15202 7039 15518 7040
rect 2245 6560 2561 6561
rect 2245 6496 2251 6560
rect 2315 6496 2331 6560
rect 2395 6496 2411 6560
rect 2475 6496 2491 6560
rect 2555 6496 2561 6560
rect 2245 6495 2561 6496
rect 5947 6560 6263 6561
rect 5947 6496 5953 6560
rect 6017 6496 6033 6560
rect 6097 6496 6113 6560
rect 6177 6496 6193 6560
rect 6257 6496 6263 6560
rect 5947 6495 6263 6496
rect 9649 6560 9965 6561
rect 9649 6496 9655 6560
rect 9719 6496 9735 6560
rect 9799 6496 9815 6560
rect 9879 6496 9895 6560
rect 9959 6496 9965 6560
rect 9649 6495 9965 6496
rect 13351 6560 13667 6561
rect 13351 6496 13357 6560
rect 13421 6496 13437 6560
rect 13501 6496 13517 6560
rect 13581 6496 13597 6560
rect 13661 6496 13667 6560
rect 13351 6495 13667 6496
rect 4096 6016 4412 6017
rect 4096 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4342 6016
rect 4406 5952 4412 6016
rect 4096 5951 4412 5952
rect 7798 6016 8114 6017
rect 7798 5952 7804 6016
rect 7868 5952 7884 6016
rect 7948 5952 7964 6016
rect 8028 5952 8044 6016
rect 8108 5952 8114 6016
rect 7798 5951 8114 5952
rect 11500 6016 11816 6017
rect 11500 5952 11506 6016
rect 11570 5952 11586 6016
rect 11650 5952 11666 6016
rect 11730 5952 11746 6016
rect 11810 5952 11816 6016
rect 11500 5951 11816 5952
rect 15202 6016 15518 6017
rect 15202 5952 15208 6016
rect 15272 5952 15288 6016
rect 15352 5952 15368 6016
rect 15432 5952 15448 6016
rect 15512 5952 15518 6016
rect 15202 5951 15518 5952
rect 2245 5472 2561 5473
rect 2245 5408 2251 5472
rect 2315 5408 2331 5472
rect 2395 5408 2411 5472
rect 2475 5408 2491 5472
rect 2555 5408 2561 5472
rect 2245 5407 2561 5408
rect 5947 5472 6263 5473
rect 5947 5408 5953 5472
rect 6017 5408 6033 5472
rect 6097 5408 6113 5472
rect 6177 5408 6193 5472
rect 6257 5408 6263 5472
rect 5947 5407 6263 5408
rect 9649 5472 9965 5473
rect 9649 5408 9655 5472
rect 9719 5408 9735 5472
rect 9799 5408 9815 5472
rect 9879 5408 9895 5472
rect 9959 5408 9965 5472
rect 9649 5407 9965 5408
rect 13351 5472 13667 5473
rect 13351 5408 13357 5472
rect 13421 5408 13437 5472
rect 13501 5408 13517 5472
rect 13581 5408 13597 5472
rect 13661 5408 13667 5472
rect 13351 5407 13667 5408
rect 4096 4928 4412 4929
rect 4096 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4342 4928
rect 4406 4864 4412 4928
rect 4096 4863 4412 4864
rect 7798 4928 8114 4929
rect 7798 4864 7804 4928
rect 7868 4864 7884 4928
rect 7948 4864 7964 4928
rect 8028 4864 8044 4928
rect 8108 4864 8114 4928
rect 7798 4863 8114 4864
rect 11500 4928 11816 4929
rect 11500 4864 11506 4928
rect 11570 4864 11586 4928
rect 11650 4864 11666 4928
rect 11730 4864 11746 4928
rect 11810 4864 11816 4928
rect 11500 4863 11816 4864
rect 15202 4928 15518 4929
rect 15202 4864 15208 4928
rect 15272 4864 15288 4928
rect 15352 4864 15368 4928
rect 15432 4864 15448 4928
rect 15512 4864 15518 4928
rect 15202 4863 15518 4864
rect 2245 4384 2561 4385
rect 2245 4320 2251 4384
rect 2315 4320 2331 4384
rect 2395 4320 2411 4384
rect 2475 4320 2491 4384
rect 2555 4320 2561 4384
rect 2245 4319 2561 4320
rect 5947 4384 6263 4385
rect 5947 4320 5953 4384
rect 6017 4320 6033 4384
rect 6097 4320 6113 4384
rect 6177 4320 6193 4384
rect 6257 4320 6263 4384
rect 5947 4319 6263 4320
rect 9649 4384 9965 4385
rect 9649 4320 9655 4384
rect 9719 4320 9735 4384
rect 9799 4320 9815 4384
rect 9879 4320 9895 4384
rect 9959 4320 9965 4384
rect 9649 4319 9965 4320
rect 13351 4384 13667 4385
rect 13351 4320 13357 4384
rect 13421 4320 13437 4384
rect 13501 4320 13517 4384
rect 13581 4320 13597 4384
rect 13661 4320 13667 4384
rect 13351 4319 13667 4320
rect 11237 4178 11303 4181
rect 11237 4176 15578 4178
rect 11237 4120 11242 4176
rect 11298 4170 15578 4176
rect 11298 4120 15946 4170
rect 11237 4118 15946 4120
rect 11237 4115 11303 4118
rect 15518 4110 15946 4118
rect 15886 3936 15946 4110
rect 4096 3840 4412 3841
rect 4096 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4342 3840
rect 4406 3776 4412 3840
rect 4096 3775 4412 3776
rect 7798 3840 8114 3841
rect 7798 3776 7804 3840
rect 7868 3776 7884 3840
rect 7948 3776 7964 3840
rect 8028 3776 8044 3840
rect 8108 3776 8114 3840
rect 7798 3775 8114 3776
rect 11500 3840 11816 3841
rect 11500 3776 11506 3840
rect 11570 3776 11586 3840
rect 11650 3776 11666 3840
rect 11730 3776 11746 3840
rect 11810 3776 11816 3840
rect 11500 3775 11816 3776
rect 15202 3840 15518 3841
rect 15202 3776 15208 3840
rect 15272 3776 15288 3840
rect 15352 3776 15368 3840
rect 15432 3776 15448 3840
rect 15512 3776 15518 3840
rect 15600 3816 16000 3936
rect 15202 3775 15518 3776
rect 2245 3296 2561 3297
rect 2245 3232 2251 3296
rect 2315 3232 2331 3296
rect 2395 3232 2411 3296
rect 2475 3232 2491 3296
rect 2555 3232 2561 3296
rect 2245 3231 2561 3232
rect 5947 3296 6263 3297
rect 5947 3232 5953 3296
rect 6017 3232 6033 3296
rect 6097 3232 6113 3296
rect 6177 3232 6193 3296
rect 6257 3232 6263 3296
rect 5947 3231 6263 3232
rect 9649 3296 9965 3297
rect 9649 3232 9655 3296
rect 9719 3232 9735 3296
rect 9799 3232 9815 3296
rect 9879 3232 9895 3296
rect 9959 3232 9965 3296
rect 9649 3231 9965 3232
rect 13351 3296 13667 3297
rect 13351 3232 13357 3296
rect 13421 3232 13437 3296
rect 13501 3232 13517 3296
rect 13581 3232 13597 3296
rect 13661 3232 13667 3296
rect 13351 3231 13667 3232
rect 4096 2752 4412 2753
rect 4096 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4342 2752
rect 4406 2688 4412 2752
rect 4096 2687 4412 2688
rect 7798 2752 8114 2753
rect 7798 2688 7804 2752
rect 7868 2688 7884 2752
rect 7948 2688 7964 2752
rect 8028 2688 8044 2752
rect 8108 2688 8114 2752
rect 7798 2687 8114 2688
rect 11500 2752 11816 2753
rect 11500 2688 11506 2752
rect 11570 2688 11586 2752
rect 11650 2688 11666 2752
rect 11730 2688 11746 2752
rect 11810 2688 11816 2752
rect 11500 2687 11816 2688
rect 15202 2752 15518 2753
rect 15202 2688 15208 2752
rect 15272 2688 15288 2752
rect 15352 2688 15368 2752
rect 15432 2688 15448 2752
rect 15512 2688 15518 2752
rect 15202 2687 15518 2688
rect 2245 2208 2561 2209
rect 2245 2144 2251 2208
rect 2315 2144 2331 2208
rect 2395 2144 2411 2208
rect 2475 2144 2491 2208
rect 2555 2144 2561 2208
rect 2245 2143 2561 2144
rect 5947 2208 6263 2209
rect 5947 2144 5953 2208
rect 6017 2144 6033 2208
rect 6097 2144 6113 2208
rect 6177 2144 6193 2208
rect 6257 2144 6263 2208
rect 5947 2143 6263 2144
rect 9649 2208 9965 2209
rect 9649 2144 9655 2208
rect 9719 2144 9735 2208
rect 9799 2144 9815 2208
rect 9879 2144 9895 2208
rect 9959 2144 9965 2208
rect 9649 2143 9965 2144
rect 13351 2208 13667 2209
rect 13351 2144 13357 2208
rect 13421 2144 13437 2208
rect 13501 2144 13517 2208
rect 13581 2144 13597 2208
rect 13661 2144 13667 2208
rect 13351 2143 13667 2144
rect 4096 1664 4412 1665
rect 4096 1600 4102 1664
rect 4166 1600 4182 1664
rect 4246 1600 4262 1664
rect 4326 1600 4342 1664
rect 4406 1600 4412 1664
rect 4096 1599 4412 1600
rect 7798 1664 8114 1665
rect 7798 1600 7804 1664
rect 7868 1600 7884 1664
rect 7948 1600 7964 1664
rect 8028 1600 8044 1664
rect 8108 1600 8114 1664
rect 7798 1599 8114 1600
rect 11500 1664 11816 1665
rect 11500 1600 11506 1664
rect 11570 1600 11586 1664
rect 11650 1600 11666 1664
rect 11730 1600 11746 1664
rect 11810 1600 11816 1664
rect 11500 1599 11816 1600
rect 15202 1664 15518 1665
rect 15202 1600 15208 1664
rect 15272 1600 15288 1664
rect 15352 1600 15368 1664
rect 15432 1600 15448 1664
rect 15512 1600 15518 1664
rect 15202 1599 15518 1600
rect 2245 1120 2561 1121
rect 2245 1056 2251 1120
rect 2315 1056 2331 1120
rect 2395 1056 2411 1120
rect 2475 1056 2491 1120
rect 2555 1056 2561 1120
rect 2245 1055 2561 1056
rect 5947 1120 6263 1121
rect 5947 1056 5953 1120
rect 6017 1056 6033 1120
rect 6097 1056 6113 1120
rect 6177 1056 6193 1120
rect 6257 1056 6263 1120
rect 5947 1055 6263 1056
rect 9649 1120 9965 1121
rect 9649 1056 9655 1120
rect 9719 1056 9735 1120
rect 9799 1056 9815 1120
rect 9879 1056 9895 1120
rect 9959 1056 9965 1120
rect 9649 1055 9965 1056
rect 13351 1120 13667 1121
rect 13351 1056 13357 1120
rect 13421 1056 13437 1120
rect 13501 1056 13517 1120
rect 13581 1056 13597 1120
rect 13661 1056 13667 1120
rect 13351 1055 13667 1056
rect 4096 576 4412 577
rect 4096 512 4102 576
rect 4166 512 4182 576
rect 4246 512 4262 576
rect 4326 512 4342 576
rect 4406 512 4412 576
rect 4096 511 4412 512
rect 7798 576 8114 577
rect 7798 512 7804 576
rect 7868 512 7884 576
rect 7948 512 7964 576
rect 8028 512 8044 576
rect 8108 512 8114 576
rect 7798 511 8114 512
rect 11500 576 11816 577
rect 11500 512 11506 576
rect 11570 512 11586 576
rect 11650 512 11666 576
rect 11730 512 11746 576
rect 11810 512 11816 576
rect 11500 511 11816 512
rect 15202 576 15518 577
rect 15202 512 15208 576
rect 15272 512 15288 576
rect 15352 512 15368 576
rect 15432 512 15448 576
rect 15512 512 15518 576
rect 15202 511 15518 512
<< via3 >>
rect 2251 15260 2315 15264
rect 2251 15204 2255 15260
rect 2255 15204 2311 15260
rect 2311 15204 2315 15260
rect 2251 15200 2315 15204
rect 2331 15260 2395 15264
rect 2331 15204 2335 15260
rect 2335 15204 2391 15260
rect 2391 15204 2395 15260
rect 2331 15200 2395 15204
rect 2411 15260 2475 15264
rect 2411 15204 2415 15260
rect 2415 15204 2471 15260
rect 2471 15204 2475 15260
rect 2411 15200 2475 15204
rect 2491 15260 2555 15264
rect 2491 15204 2495 15260
rect 2495 15204 2551 15260
rect 2551 15204 2555 15260
rect 2491 15200 2555 15204
rect 5953 15260 6017 15264
rect 5953 15204 5957 15260
rect 5957 15204 6013 15260
rect 6013 15204 6017 15260
rect 5953 15200 6017 15204
rect 6033 15260 6097 15264
rect 6033 15204 6037 15260
rect 6037 15204 6093 15260
rect 6093 15204 6097 15260
rect 6033 15200 6097 15204
rect 6113 15260 6177 15264
rect 6113 15204 6117 15260
rect 6117 15204 6173 15260
rect 6173 15204 6177 15260
rect 6113 15200 6177 15204
rect 6193 15260 6257 15264
rect 6193 15204 6197 15260
rect 6197 15204 6253 15260
rect 6253 15204 6257 15260
rect 6193 15200 6257 15204
rect 9655 15260 9719 15264
rect 9655 15204 9659 15260
rect 9659 15204 9715 15260
rect 9715 15204 9719 15260
rect 9655 15200 9719 15204
rect 9735 15260 9799 15264
rect 9735 15204 9739 15260
rect 9739 15204 9795 15260
rect 9795 15204 9799 15260
rect 9735 15200 9799 15204
rect 9815 15260 9879 15264
rect 9815 15204 9819 15260
rect 9819 15204 9875 15260
rect 9875 15204 9879 15260
rect 9815 15200 9879 15204
rect 9895 15260 9959 15264
rect 9895 15204 9899 15260
rect 9899 15204 9955 15260
rect 9955 15204 9959 15260
rect 9895 15200 9959 15204
rect 13357 15260 13421 15264
rect 13357 15204 13361 15260
rect 13361 15204 13417 15260
rect 13417 15204 13421 15260
rect 13357 15200 13421 15204
rect 13437 15260 13501 15264
rect 13437 15204 13441 15260
rect 13441 15204 13497 15260
rect 13497 15204 13501 15260
rect 13437 15200 13501 15204
rect 13517 15260 13581 15264
rect 13517 15204 13521 15260
rect 13521 15204 13577 15260
rect 13577 15204 13581 15260
rect 13517 15200 13581 15204
rect 13597 15260 13661 15264
rect 13597 15204 13601 15260
rect 13601 15204 13657 15260
rect 13657 15204 13661 15260
rect 13597 15200 13661 15204
rect 4102 14716 4166 14720
rect 4102 14660 4106 14716
rect 4106 14660 4162 14716
rect 4162 14660 4166 14716
rect 4102 14656 4166 14660
rect 4182 14716 4246 14720
rect 4182 14660 4186 14716
rect 4186 14660 4242 14716
rect 4242 14660 4246 14716
rect 4182 14656 4246 14660
rect 4262 14716 4326 14720
rect 4262 14660 4266 14716
rect 4266 14660 4322 14716
rect 4322 14660 4326 14716
rect 4262 14656 4326 14660
rect 4342 14716 4406 14720
rect 4342 14660 4346 14716
rect 4346 14660 4402 14716
rect 4402 14660 4406 14716
rect 4342 14656 4406 14660
rect 7804 14716 7868 14720
rect 7804 14660 7808 14716
rect 7808 14660 7864 14716
rect 7864 14660 7868 14716
rect 7804 14656 7868 14660
rect 7884 14716 7948 14720
rect 7884 14660 7888 14716
rect 7888 14660 7944 14716
rect 7944 14660 7948 14716
rect 7884 14656 7948 14660
rect 7964 14716 8028 14720
rect 7964 14660 7968 14716
rect 7968 14660 8024 14716
rect 8024 14660 8028 14716
rect 7964 14656 8028 14660
rect 8044 14716 8108 14720
rect 8044 14660 8048 14716
rect 8048 14660 8104 14716
rect 8104 14660 8108 14716
rect 8044 14656 8108 14660
rect 11506 14716 11570 14720
rect 11506 14660 11510 14716
rect 11510 14660 11566 14716
rect 11566 14660 11570 14716
rect 11506 14656 11570 14660
rect 11586 14716 11650 14720
rect 11586 14660 11590 14716
rect 11590 14660 11646 14716
rect 11646 14660 11650 14716
rect 11586 14656 11650 14660
rect 11666 14716 11730 14720
rect 11666 14660 11670 14716
rect 11670 14660 11726 14716
rect 11726 14660 11730 14716
rect 11666 14656 11730 14660
rect 11746 14716 11810 14720
rect 11746 14660 11750 14716
rect 11750 14660 11806 14716
rect 11806 14660 11810 14716
rect 11746 14656 11810 14660
rect 15208 14716 15272 14720
rect 15208 14660 15212 14716
rect 15212 14660 15268 14716
rect 15268 14660 15272 14716
rect 15208 14656 15272 14660
rect 15288 14716 15352 14720
rect 15288 14660 15292 14716
rect 15292 14660 15348 14716
rect 15348 14660 15352 14716
rect 15288 14656 15352 14660
rect 15368 14716 15432 14720
rect 15368 14660 15372 14716
rect 15372 14660 15428 14716
rect 15428 14660 15432 14716
rect 15368 14656 15432 14660
rect 15448 14716 15512 14720
rect 15448 14660 15452 14716
rect 15452 14660 15508 14716
rect 15508 14660 15512 14716
rect 15448 14656 15512 14660
rect 2251 14172 2315 14176
rect 2251 14116 2255 14172
rect 2255 14116 2311 14172
rect 2311 14116 2315 14172
rect 2251 14112 2315 14116
rect 2331 14172 2395 14176
rect 2331 14116 2335 14172
rect 2335 14116 2391 14172
rect 2391 14116 2395 14172
rect 2331 14112 2395 14116
rect 2411 14172 2475 14176
rect 2411 14116 2415 14172
rect 2415 14116 2471 14172
rect 2471 14116 2475 14172
rect 2411 14112 2475 14116
rect 2491 14172 2555 14176
rect 2491 14116 2495 14172
rect 2495 14116 2551 14172
rect 2551 14116 2555 14172
rect 2491 14112 2555 14116
rect 5953 14172 6017 14176
rect 5953 14116 5957 14172
rect 5957 14116 6013 14172
rect 6013 14116 6017 14172
rect 5953 14112 6017 14116
rect 6033 14172 6097 14176
rect 6033 14116 6037 14172
rect 6037 14116 6093 14172
rect 6093 14116 6097 14172
rect 6033 14112 6097 14116
rect 6113 14172 6177 14176
rect 6113 14116 6117 14172
rect 6117 14116 6173 14172
rect 6173 14116 6177 14172
rect 6113 14112 6177 14116
rect 6193 14172 6257 14176
rect 6193 14116 6197 14172
rect 6197 14116 6253 14172
rect 6253 14116 6257 14172
rect 6193 14112 6257 14116
rect 9655 14172 9719 14176
rect 9655 14116 9659 14172
rect 9659 14116 9715 14172
rect 9715 14116 9719 14172
rect 9655 14112 9719 14116
rect 9735 14172 9799 14176
rect 9735 14116 9739 14172
rect 9739 14116 9795 14172
rect 9795 14116 9799 14172
rect 9735 14112 9799 14116
rect 9815 14172 9879 14176
rect 9815 14116 9819 14172
rect 9819 14116 9875 14172
rect 9875 14116 9879 14172
rect 9815 14112 9879 14116
rect 9895 14172 9959 14176
rect 9895 14116 9899 14172
rect 9899 14116 9955 14172
rect 9955 14116 9959 14172
rect 9895 14112 9959 14116
rect 13357 14172 13421 14176
rect 13357 14116 13361 14172
rect 13361 14116 13417 14172
rect 13417 14116 13421 14172
rect 13357 14112 13421 14116
rect 13437 14172 13501 14176
rect 13437 14116 13441 14172
rect 13441 14116 13497 14172
rect 13497 14116 13501 14172
rect 13437 14112 13501 14116
rect 13517 14172 13581 14176
rect 13517 14116 13521 14172
rect 13521 14116 13577 14172
rect 13577 14116 13581 14172
rect 13517 14112 13581 14116
rect 13597 14172 13661 14176
rect 13597 14116 13601 14172
rect 13601 14116 13657 14172
rect 13657 14116 13661 14172
rect 13597 14112 13661 14116
rect 4102 13628 4166 13632
rect 4102 13572 4106 13628
rect 4106 13572 4162 13628
rect 4162 13572 4166 13628
rect 4102 13568 4166 13572
rect 4182 13628 4246 13632
rect 4182 13572 4186 13628
rect 4186 13572 4242 13628
rect 4242 13572 4246 13628
rect 4182 13568 4246 13572
rect 4262 13628 4326 13632
rect 4262 13572 4266 13628
rect 4266 13572 4322 13628
rect 4322 13572 4326 13628
rect 4262 13568 4326 13572
rect 4342 13628 4406 13632
rect 4342 13572 4346 13628
rect 4346 13572 4402 13628
rect 4402 13572 4406 13628
rect 4342 13568 4406 13572
rect 7804 13628 7868 13632
rect 7804 13572 7808 13628
rect 7808 13572 7864 13628
rect 7864 13572 7868 13628
rect 7804 13568 7868 13572
rect 7884 13628 7948 13632
rect 7884 13572 7888 13628
rect 7888 13572 7944 13628
rect 7944 13572 7948 13628
rect 7884 13568 7948 13572
rect 7964 13628 8028 13632
rect 7964 13572 7968 13628
rect 7968 13572 8024 13628
rect 8024 13572 8028 13628
rect 7964 13568 8028 13572
rect 8044 13628 8108 13632
rect 8044 13572 8048 13628
rect 8048 13572 8104 13628
rect 8104 13572 8108 13628
rect 8044 13568 8108 13572
rect 11506 13628 11570 13632
rect 11506 13572 11510 13628
rect 11510 13572 11566 13628
rect 11566 13572 11570 13628
rect 11506 13568 11570 13572
rect 11586 13628 11650 13632
rect 11586 13572 11590 13628
rect 11590 13572 11646 13628
rect 11646 13572 11650 13628
rect 11586 13568 11650 13572
rect 11666 13628 11730 13632
rect 11666 13572 11670 13628
rect 11670 13572 11726 13628
rect 11726 13572 11730 13628
rect 11666 13568 11730 13572
rect 11746 13628 11810 13632
rect 11746 13572 11750 13628
rect 11750 13572 11806 13628
rect 11806 13572 11810 13628
rect 11746 13568 11810 13572
rect 15208 13628 15272 13632
rect 15208 13572 15212 13628
rect 15212 13572 15268 13628
rect 15268 13572 15272 13628
rect 15208 13568 15272 13572
rect 15288 13628 15352 13632
rect 15288 13572 15292 13628
rect 15292 13572 15348 13628
rect 15348 13572 15352 13628
rect 15288 13568 15352 13572
rect 15368 13628 15432 13632
rect 15368 13572 15372 13628
rect 15372 13572 15428 13628
rect 15428 13572 15432 13628
rect 15368 13568 15432 13572
rect 15448 13628 15512 13632
rect 15448 13572 15452 13628
rect 15452 13572 15508 13628
rect 15508 13572 15512 13628
rect 15448 13568 15512 13572
rect 2251 13084 2315 13088
rect 2251 13028 2255 13084
rect 2255 13028 2311 13084
rect 2311 13028 2315 13084
rect 2251 13024 2315 13028
rect 2331 13084 2395 13088
rect 2331 13028 2335 13084
rect 2335 13028 2391 13084
rect 2391 13028 2395 13084
rect 2331 13024 2395 13028
rect 2411 13084 2475 13088
rect 2411 13028 2415 13084
rect 2415 13028 2471 13084
rect 2471 13028 2475 13084
rect 2411 13024 2475 13028
rect 2491 13084 2555 13088
rect 2491 13028 2495 13084
rect 2495 13028 2551 13084
rect 2551 13028 2555 13084
rect 2491 13024 2555 13028
rect 5953 13084 6017 13088
rect 5953 13028 5957 13084
rect 5957 13028 6013 13084
rect 6013 13028 6017 13084
rect 5953 13024 6017 13028
rect 6033 13084 6097 13088
rect 6033 13028 6037 13084
rect 6037 13028 6093 13084
rect 6093 13028 6097 13084
rect 6033 13024 6097 13028
rect 6113 13084 6177 13088
rect 6113 13028 6117 13084
rect 6117 13028 6173 13084
rect 6173 13028 6177 13084
rect 6113 13024 6177 13028
rect 6193 13084 6257 13088
rect 6193 13028 6197 13084
rect 6197 13028 6253 13084
rect 6253 13028 6257 13084
rect 6193 13024 6257 13028
rect 9655 13084 9719 13088
rect 9655 13028 9659 13084
rect 9659 13028 9715 13084
rect 9715 13028 9719 13084
rect 9655 13024 9719 13028
rect 9735 13084 9799 13088
rect 9735 13028 9739 13084
rect 9739 13028 9795 13084
rect 9795 13028 9799 13084
rect 9735 13024 9799 13028
rect 9815 13084 9879 13088
rect 9815 13028 9819 13084
rect 9819 13028 9875 13084
rect 9875 13028 9879 13084
rect 9815 13024 9879 13028
rect 9895 13084 9959 13088
rect 9895 13028 9899 13084
rect 9899 13028 9955 13084
rect 9955 13028 9959 13084
rect 9895 13024 9959 13028
rect 13357 13084 13421 13088
rect 13357 13028 13361 13084
rect 13361 13028 13417 13084
rect 13417 13028 13421 13084
rect 13357 13024 13421 13028
rect 13437 13084 13501 13088
rect 13437 13028 13441 13084
rect 13441 13028 13497 13084
rect 13497 13028 13501 13084
rect 13437 13024 13501 13028
rect 13517 13084 13581 13088
rect 13517 13028 13521 13084
rect 13521 13028 13577 13084
rect 13577 13028 13581 13084
rect 13517 13024 13581 13028
rect 13597 13084 13661 13088
rect 13597 13028 13601 13084
rect 13601 13028 13657 13084
rect 13657 13028 13661 13084
rect 13597 13024 13661 13028
rect 4102 12540 4166 12544
rect 4102 12484 4106 12540
rect 4106 12484 4162 12540
rect 4162 12484 4166 12540
rect 4102 12480 4166 12484
rect 4182 12540 4246 12544
rect 4182 12484 4186 12540
rect 4186 12484 4242 12540
rect 4242 12484 4246 12540
rect 4182 12480 4246 12484
rect 4262 12540 4326 12544
rect 4262 12484 4266 12540
rect 4266 12484 4322 12540
rect 4322 12484 4326 12540
rect 4262 12480 4326 12484
rect 4342 12540 4406 12544
rect 4342 12484 4346 12540
rect 4346 12484 4402 12540
rect 4402 12484 4406 12540
rect 4342 12480 4406 12484
rect 7804 12540 7868 12544
rect 7804 12484 7808 12540
rect 7808 12484 7864 12540
rect 7864 12484 7868 12540
rect 7804 12480 7868 12484
rect 7884 12540 7948 12544
rect 7884 12484 7888 12540
rect 7888 12484 7944 12540
rect 7944 12484 7948 12540
rect 7884 12480 7948 12484
rect 7964 12540 8028 12544
rect 7964 12484 7968 12540
rect 7968 12484 8024 12540
rect 8024 12484 8028 12540
rect 7964 12480 8028 12484
rect 8044 12540 8108 12544
rect 8044 12484 8048 12540
rect 8048 12484 8104 12540
rect 8104 12484 8108 12540
rect 8044 12480 8108 12484
rect 11506 12540 11570 12544
rect 11506 12484 11510 12540
rect 11510 12484 11566 12540
rect 11566 12484 11570 12540
rect 11506 12480 11570 12484
rect 11586 12540 11650 12544
rect 11586 12484 11590 12540
rect 11590 12484 11646 12540
rect 11646 12484 11650 12540
rect 11586 12480 11650 12484
rect 11666 12540 11730 12544
rect 11666 12484 11670 12540
rect 11670 12484 11726 12540
rect 11726 12484 11730 12540
rect 11666 12480 11730 12484
rect 11746 12540 11810 12544
rect 11746 12484 11750 12540
rect 11750 12484 11806 12540
rect 11806 12484 11810 12540
rect 11746 12480 11810 12484
rect 15208 12540 15272 12544
rect 15208 12484 15212 12540
rect 15212 12484 15268 12540
rect 15268 12484 15272 12540
rect 15208 12480 15272 12484
rect 15288 12540 15352 12544
rect 15288 12484 15292 12540
rect 15292 12484 15348 12540
rect 15348 12484 15352 12540
rect 15288 12480 15352 12484
rect 15368 12540 15432 12544
rect 15368 12484 15372 12540
rect 15372 12484 15428 12540
rect 15428 12484 15432 12540
rect 15368 12480 15432 12484
rect 15448 12540 15512 12544
rect 15448 12484 15452 12540
rect 15452 12484 15508 12540
rect 15508 12484 15512 12540
rect 15448 12480 15512 12484
rect 2251 11996 2315 12000
rect 2251 11940 2255 11996
rect 2255 11940 2311 11996
rect 2311 11940 2315 11996
rect 2251 11936 2315 11940
rect 2331 11996 2395 12000
rect 2331 11940 2335 11996
rect 2335 11940 2391 11996
rect 2391 11940 2395 11996
rect 2331 11936 2395 11940
rect 2411 11996 2475 12000
rect 2411 11940 2415 11996
rect 2415 11940 2471 11996
rect 2471 11940 2475 11996
rect 2411 11936 2475 11940
rect 2491 11996 2555 12000
rect 2491 11940 2495 11996
rect 2495 11940 2551 11996
rect 2551 11940 2555 11996
rect 2491 11936 2555 11940
rect 5953 11996 6017 12000
rect 5953 11940 5957 11996
rect 5957 11940 6013 11996
rect 6013 11940 6017 11996
rect 5953 11936 6017 11940
rect 6033 11996 6097 12000
rect 6033 11940 6037 11996
rect 6037 11940 6093 11996
rect 6093 11940 6097 11996
rect 6033 11936 6097 11940
rect 6113 11996 6177 12000
rect 6113 11940 6117 11996
rect 6117 11940 6173 11996
rect 6173 11940 6177 11996
rect 6113 11936 6177 11940
rect 6193 11996 6257 12000
rect 6193 11940 6197 11996
rect 6197 11940 6253 11996
rect 6253 11940 6257 11996
rect 6193 11936 6257 11940
rect 9655 11996 9719 12000
rect 9655 11940 9659 11996
rect 9659 11940 9715 11996
rect 9715 11940 9719 11996
rect 9655 11936 9719 11940
rect 9735 11996 9799 12000
rect 9735 11940 9739 11996
rect 9739 11940 9795 11996
rect 9795 11940 9799 11996
rect 9735 11936 9799 11940
rect 9815 11996 9879 12000
rect 9815 11940 9819 11996
rect 9819 11940 9875 11996
rect 9875 11940 9879 11996
rect 9815 11936 9879 11940
rect 9895 11996 9959 12000
rect 9895 11940 9899 11996
rect 9899 11940 9955 11996
rect 9955 11940 9959 11996
rect 9895 11936 9959 11940
rect 13357 11996 13421 12000
rect 13357 11940 13361 11996
rect 13361 11940 13417 11996
rect 13417 11940 13421 11996
rect 13357 11936 13421 11940
rect 13437 11996 13501 12000
rect 13437 11940 13441 11996
rect 13441 11940 13497 11996
rect 13497 11940 13501 11996
rect 13437 11936 13501 11940
rect 13517 11996 13581 12000
rect 13517 11940 13521 11996
rect 13521 11940 13577 11996
rect 13577 11940 13581 11996
rect 13517 11936 13581 11940
rect 13597 11996 13661 12000
rect 13597 11940 13601 11996
rect 13601 11940 13657 11996
rect 13657 11940 13661 11996
rect 13597 11936 13661 11940
rect 4102 11452 4166 11456
rect 4102 11396 4106 11452
rect 4106 11396 4162 11452
rect 4162 11396 4166 11452
rect 4102 11392 4166 11396
rect 4182 11452 4246 11456
rect 4182 11396 4186 11452
rect 4186 11396 4242 11452
rect 4242 11396 4246 11452
rect 4182 11392 4246 11396
rect 4262 11452 4326 11456
rect 4262 11396 4266 11452
rect 4266 11396 4322 11452
rect 4322 11396 4326 11452
rect 4262 11392 4326 11396
rect 4342 11452 4406 11456
rect 4342 11396 4346 11452
rect 4346 11396 4402 11452
rect 4402 11396 4406 11452
rect 4342 11392 4406 11396
rect 7804 11452 7868 11456
rect 7804 11396 7808 11452
rect 7808 11396 7864 11452
rect 7864 11396 7868 11452
rect 7804 11392 7868 11396
rect 7884 11452 7948 11456
rect 7884 11396 7888 11452
rect 7888 11396 7944 11452
rect 7944 11396 7948 11452
rect 7884 11392 7948 11396
rect 7964 11452 8028 11456
rect 7964 11396 7968 11452
rect 7968 11396 8024 11452
rect 8024 11396 8028 11452
rect 7964 11392 8028 11396
rect 8044 11452 8108 11456
rect 8044 11396 8048 11452
rect 8048 11396 8104 11452
rect 8104 11396 8108 11452
rect 8044 11392 8108 11396
rect 11506 11452 11570 11456
rect 11506 11396 11510 11452
rect 11510 11396 11566 11452
rect 11566 11396 11570 11452
rect 11506 11392 11570 11396
rect 11586 11452 11650 11456
rect 11586 11396 11590 11452
rect 11590 11396 11646 11452
rect 11646 11396 11650 11452
rect 11586 11392 11650 11396
rect 11666 11452 11730 11456
rect 11666 11396 11670 11452
rect 11670 11396 11726 11452
rect 11726 11396 11730 11452
rect 11666 11392 11730 11396
rect 11746 11452 11810 11456
rect 11746 11396 11750 11452
rect 11750 11396 11806 11452
rect 11806 11396 11810 11452
rect 11746 11392 11810 11396
rect 15208 11452 15272 11456
rect 15208 11396 15212 11452
rect 15212 11396 15268 11452
rect 15268 11396 15272 11452
rect 15208 11392 15272 11396
rect 15288 11452 15352 11456
rect 15288 11396 15292 11452
rect 15292 11396 15348 11452
rect 15348 11396 15352 11452
rect 15288 11392 15352 11396
rect 15368 11452 15432 11456
rect 15368 11396 15372 11452
rect 15372 11396 15428 11452
rect 15428 11396 15432 11452
rect 15368 11392 15432 11396
rect 15448 11452 15512 11456
rect 15448 11396 15452 11452
rect 15452 11396 15508 11452
rect 15508 11396 15512 11452
rect 15448 11392 15512 11396
rect 2251 10908 2315 10912
rect 2251 10852 2255 10908
rect 2255 10852 2311 10908
rect 2311 10852 2315 10908
rect 2251 10848 2315 10852
rect 2331 10908 2395 10912
rect 2331 10852 2335 10908
rect 2335 10852 2391 10908
rect 2391 10852 2395 10908
rect 2331 10848 2395 10852
rect 2411 10908 2475 10912
rect 2411 10852 2415 10908
rect 2415 10852 2471 10908
rect 2471 10852 2475 10908
rect 2411 10848 2475 10852
rect 2491 10908 2555 10912
rect 2491 10852 2495 10908
rect 2495 10852 2551 10908
rect 2551 10852 2555 10908
rect 2491 10848 2555 10852
rect 5953 10908 6017 10912
rect 5953 10852 5957 10908
rect 5957 10852 6013 10908
rect 6013 10852 6017 10908
rect 5953 10848 6017 10852
rect 6033 10908 6097 10912
rect 6033 10852 6037 10908
rect 6037 10852 6093 10908
rect 6093 10852 6097 10908
rect 6033 10848 6097 10852
rect 6113 10908 6177 10912
rect 6113 10852 6117 10908
rect 6117 10852 6173 10908
rect 6173 10852 6177 10908
rect 6113 10848 6177 10852
rect 6193 10908 6257 10912
rect 6193 10852 6197 10908
rect 6197 10852 6253 10908
rect 6253 10852 6257 10908
rect 6193 10848 6257 10852
rect 9655 10908 9719 10912
rect 9655 10852 9659 10908
rect 9659 10852 9715 10908
rect 9715 10852 9719 10908
rect 9655 10848 9719 10852
rect 9735 10908 9799 10912
rect 9735 10852 9739 10908
rect 9739 10852 9795 10908
rect 9795 10852 9799 10908
rect 9735 10848 9799 10852
rect 9815 10908 9879 10912
rect 9815 10852 9819 10908
rect 9819 10852 9875 10908
rect 9875 10852 9879 10908
rect 9815 10848 9879 10852
rect 9895 10908 9959 10912
rect 9895 10852 9899 10908
rect 9899 10852 9955 10908
rect 9955 10852 9959 10908
rect 9895 10848 9959 10852
rect 13357 10908 13421 10912
rect 13357 10852 13361 10908
rect 13361 10852 13417 10908
rect 13417 10852 13421 10908
rect 13357 10848 13421 10852
rect 13437 10908 13501 10912
rect 13437 10852 13441 10908
rect 13441 10852 13497 10908
rect 13497 10852 13501 10908
rect 13437 10848 13501 10852
rect 13517 10908 13581 10912
rect 13517 10852 13521 10908
rect 13521 10852 13577 10908
rect 13577 10852 13581 10908
rect 13517 10848 13581 10852
rect 13597 10908 13661 10912
rect 13597 10852 13601 10908
rect 13601 10852 13657 10908
rect 13657 10852 13661 10908
rect 13597 10848 13661 10852
rect 4102 10364 4166 10368
rect 4102 10308 4106 10364
rect 4106 10308 4162 10364
rect 4162 10308 4166 10364
rect 4102 10304 4166 10308
rect 4182 10364 4246 10368
rect 4182 10308 4186 10364
rect 4186 10308 4242 10364
rect 4242 10308 4246 10364
rect 4182 10304 4246 10308
rect 4262 10364 4326 10368
rect 4262 10308 4266 10364
rect 4266 10308 4322 10364
rect 4322 10308 4326 10364
rect 4262 10304 4326 10308
rect 4342 10364 4406 10368
rect 4342 10308 4346 10364
rect 4346 10308 4402 10364
rect 4402 10308 4406 10364
rect 4342 10304 4406 10308
rect 7804 10364 7868 10368
rect 7804 10308 7808 10364
rect 7808 10308 7864 10364
rect 7864 10308 7868 10364
rect 7804 10304 7868 10308
rect 7884 10364 7948 10368
rect 7884 10308 7888 10364
rect 7888 10308 7944 10364
rect 7944 10308 7948 10364
rect 7884 10304 7948 10308
rect 7964 10364 8028 10368
rect 7964 10308 7968 10364
rect 7968 10308 8024 10364
rect 8024 10308 8028 10364
rect 7964 10304 8028 10308
rect 8044 10364 8108 10368
rect 8044 10308 8048 10364
rect 8048 10308 8104 10364
rect 8104 10308 8108 10364
rect 8044 10304 8108 10308
rect 11506 10364 11570 10368
rect 11506 10308 11510 10364
rect 11510 10308 11566 10364
rect 11566 10308 11570 10364
rect 11506 10304 11570 10308
rect 11586 10364 11650 10368
rect 11586 10308 11590 10364
rect 11590 10308 11646 10364
rect 11646 10308 11650 10364
rect 11586 10304 11650 10308
rect 11666 10364 11730 10368
rect 11666 10308 11670 10364
rect 11670 10308 11726 10364
rect 11726 10308 11730 10364
rect 11666 10304 11730 10308
rect 11746 10364 11810 10368
rect 11746 10308 11750 10364
rect 11750 10308 11806 10364
rect 11806 10308 11810 10364
rect 11746 10304 11810 10308
rect 15208 10364 15272 10368
rect 15208 10308 15212 10364
rect 15212 10308 15268 10364
rect 15268 10308 15272 10364
rect 15208 10304 15272 10308
rect 15288 10364 15352 10368
rect 15288 10308 15292 10364
rect 15292 10308 15348 10364
rect 15348 10308 15352 10364
rect 15288 10304 15352 10308
rect 15368 10364 15432 10368
rect 15368 10308 15372 10364
rect 15372 10308 15428 10364
rect 15428 10308 15432 10364
rect 15368 10304 15432 10308
rect 15448 10364 15512 10368
rect 15448 10308 15452 10364
rect 15452 10308 15508 10364
rect 15508 10308 15512 10364
rect 15448 10304 15512 10308
rect 2251 9820 2315 9824
rect 2251 9764 2255 9820
rect 2255 9764 2311 9820
rect 2311 9764 2315 9820
rect 2251 9760 2315 9764
rect 2331 9820 2395 9824
rect 2331 9764 2335 9820
rect 2335 9764 2391 9820
rect 2391 9764 2395 9820
rect 2331 9760 2395 9764
rect 2411 9820 2475 9824
rect 2411 9764 2415 9820
rect 2415 9764 2471 9820
rect 2471 9764 2475 9820
rect 2411 9760 2475 9764
rect 2491 9820 2555 9824
rect 2491 9764 2495 9820
rect 2495 9764 2551 9820
rect 2551 9764 2555 9820
rect 2491 9760 2555 9764
rect 5953 9820 6017 9824
rect 5953 9764 5957 9820
rect 5957 9764 6013 9820
rect 6013 9764 6017 9820
rect 5953 9760 6017 9764
rect 6033 9820 6097 9824
rect 6033 9764 6037 9820
rect 6037 9764 6093 9820
rect 6093 9764 6097 9820
rect 6033 9760 6097 9764
rect 6113 9820 6177 9824
rect 6113 9764 6117 9820
rect 6117 9764 6173 9820
rect 6173 9764 6177 9820
rect 6113 9760 6177 9764
rect 6193 9820 6257 9824
rect 6193 9764 6197 9820
rect 6197 9764 6253 9820
rect 6253 9764 6257 9820
rect 6193 9760 6257 9764
rect 9655 9820 9719 9824
rect 9655 9764 9659 9820
rect 9659 9764 9715 9820
rect 9715 9764 9719 9820
rect 9655 9760 9719 9764
rect 9735 9820 9799 9824
rect 9735 9764 9739 9820
rect 9739 9764 9795 9820
rect 9795 9764 9799 9820
rect 9735 9760 9799 9764
rect 9815 9820 9879 9824
rect 9815 9764 9819 9820
rect 9819 9764 9875 9820
rect 9875 9764 9879 9820
rect 9815 9760 9879 9764
rect 9895 9820 9959 9824
rect 9895 9764 9899 9820
rect 9899 9764 9955 9820
rect 9955 9764 9959 9820
rect 9895 9760 9959 9764
rect 13357 9820 13421 9824
rect 13357 9764 13361 9820
rect 13361 9764 13417 9820
rect 13417 9764 13421 9820
rect 13357 9760 13421 9764
rect 13437 9820 13501 9824
rect 13437 9764 13441 9820
rect 13441 9764 13497 9820
rect 13497 9764 13501 9820
rect 13437 9760 13501 9764
rect 13517 9820 13581 9824
rect 13517 9764 13521 9820
rect 13521 9764 13577 9820
rect 13577 9764 13581 9820
rect 13517 9760 13581 9764
rect 13597 9820 13661 9824
rect 13597 9764 13601 9820
rect 13601 9764 13657 9820
rect 13657 9764 13661 9820
rect 13597 9760 13661 9764
rect 4102 9276 4166 9280
rect 4102 9220 4106 9276
rect 4106 9220 4162 9276
rect 4162 9220 4166 9276
rect 4102 9216 4166 9220
rect 4182 9276 4246 9280
rect 4182 9220 4186 9276
rect 4186 9220 4242 9276
rect 4242 9220 4246 9276
rect 4182 9216 4246 9220
rect 4262 9276 4326 9280
rect 4262 9220 4266 9276
rect 4266 9220 4322 9276
rect 4322 9220 4326 9276
rect 4262 9216 4326 9220
rect 4342 9276 4406 9280
rect 4342 9220 4346 9276
rect 4346 9220 4402 9276
rect 4402 9220 4406 9276
rect 4342 9216 4406 9220
rect 7804 9276 7868 9280
rect 7804 9220 7808 9276
rect 7808 9220 7864 9276
rect 7864 9220 7868 9276
rect 7804 9216 7868 9220
rect 7884 9276 7948 9280
rect 7884 9220 7888 9276
rect 7888 9220 7944 9276
rect 7944 9220 7948 9276
rect 7884 9216 7948 9220
rect 7964 9276 8028 9280
rect 7964 9220 7968 9276
rect 7968 9220 8024 9276
rect 8024 9220 8028 9276
rect 7964 9216 8028 9220
rect 8044 9276 8108 9280
rect 8044 9220 8048 9276
rect 8048 9220 8104 9276
rect 8104 9220 8108 9276
rect 8044 9216 8108 9220
rect 11506 9276 11570 9280
rect 11506 9220 11510 9276
rect 11510 9220 11566 9276
rect 11566 9220 11570 9276
rect 11506 9216 11570 9220
rect 11586 9276 11650 9280
rect 11586 9220 11590 9276
rect 11590 9220 11646 9276
rect 11646 9220 11650 9276
rect 11586 9216 11650 9220
rect 11666 9276 11730 9280
rect 11666 9220 11670 9276
rect 11670 9220 11726 9276
rect 11726 9220 11730 9276
rect 11666 9216 11730 9220
rect 11746 9276 11810 9280
rect 11746 9220 11750 9276
rect 11750 9220 11806 9276
rect 11806 9220 11810 9276
rect 11746 9216 11810 9220
rect 15208 9276 15272 9280
rect 15208 9220 15212 9276
rect 15212 9220 15268 9276
rect 15268 9220 15272 9276
rect 15208 9216 15272 9220
rect 15288 9276 15352 9280
rect 15288 9220 15292 9276
rect 15292 9220 15348 9276
rect 15348 9220 15352 9276
rect 15288 9216 15352 9220
rect 15368 9276 15432 9280
rect 15368 9220 15372 9276
rect 15372 9220 15428 9276
rect 15428 9220 15432 9276
rect 15368 9216 15432 9220
rect 15448 9276 15512 9280
rect 15448 9220 15452 9276
rect 15452 9220 15508 9276
rect 15508 9220 15512 9276
rect 15448 9216 15512 9220
rect 2251 8732 2315 8736
rect 2251 8676 2255 8732
rect 2255 8676 2311 8732
rect 2311 8676 2315 8732
rect 2251 8672 2315 8676
rect 2331 8732 2395 8736
rect 2331 8676 2335 8732
rect 2335 8676 2391 8732
rect 2391 8676 2395 8732
rect 2331 8672 2395 8676
rect 2411 8732 2475 8736
rect 2411 8676 2415 8732
rect 2415 8676 2471 8732
rect 2471 8676 2475 8732
rect 2411 8672 2475 8676
rect 2491 8732 2555 8736
rect 2491 8676 2495 8732
rect 2495 8676 2551 8732
rect 2551 8676 2555 8732
rect 2491 8672 2555 8676
rect 5953 8732 6017 8736
rect 5953 8676 5957 8732
rect 5957 8676 6013 8732
rect 6013 8676 6017 8732
rect 5953 8672 6017 8676
rect 6033 8732 6097 8736
rect 6033 8676 6037 8732
rect 6037 8676 6093 8732
rect 6093 8676 6097 8732
rect 6033 8672 6097 8676
rect 6113 8732 6177 8736
rect 6113 8676 6117 8732
rect 6117 8676 6173 8732
rect 6173 8676 6177 8732
rect 6113 8672 6177 8676
rect 6193 8732 6257 8736
rect 6193 8676 6197 8732
rect 6197 8676 6253 8732
rect 6253 8676 6257 8732
rect 6193 8672 6257 8676
rect 9655 8732 9719 8736
rect 9655 8676 9659 8732
rect 9659 8676 9715 8732
rect 9715 8676 9719 8732
rect 9655 8672 9719 8676
rect 9735 8732 9799 8736
rect 9735 8676 9739 8732
rect 9739 8676 9795 8732
rect 9795 8676 9799 8732
rect 9735 8672 9799 8676
rect 9815 8732 9879 8736
rect 9815 8676 9819 8732
rect 9819 8676 9875 8732
rect 9875 8676 9879 8732
rect 9815 8672 9879 8676
rect 9895 8732 9959 8736
rect 9895 8676 9899 8732
rect 9899 8676 9955 8732
rect 9955 8676 9959 8732
rect 9895 8672 9959 8676
rect 13357 8732 13421 8736
rect 13357 8676 13361 8732
rect 13361 8676 13417 8732
rect 13417 8676 13421 8732
rect 13357 8672 13421 8676
rect 13437 8732 13501 8736
rect 13437 8676 13441 8732
rect 13441 8676 13497 8732
rect 13497 8676 13501 8732
rect 13437 8672 13501 8676
rect 13517 8732 13581 8736
rect 13517 8676 13521 8732
rect 13521 8676 13577 8732
rect 13577 8676 13581 8732
rect 13517 8672 13581 8676
rect 13597 8732 13661 8736
rect 13597 8676 13601 8732
rect 13601 8676 13657 8732
rect 13657 8676 13661 8732
rect 13597 8672 13661 8676
rect 4102 8188 4166 8192
rect 4102 8132 4106 8188
rect 4106 8132 4162 8188
rect 4162 8132 4166 8188
rect 4102 8128 4166 8132
rect 4182 8188 4246 8192
rect 4182 8132 4186 8188
rect 4186 8132 4242 8188
rect 4242 8132 4246 8188
rect 4182 8128 4246 8132
rect 4262 8188 4326 8192
rect 4262 8132 4266 8188
rect 4266 8132 4322 8188
rect 4322 8132 4326 8188
rect 4262 8128 4326 8132
rect 4342 8188 4406 8192
rect 4342 8132 4346 8188
rect 4346 8132 4402 8188
rect 4402 8132 4406 8188
rect 4342 8128 4406 8132
rect 7804 8188 7868 8192
rect 7804 8132 7808 8188
rect 7808 8132 7864 8188
rect 7864 8132 7868 8188
rect 7804 8128 7868 8132
rect 7884 8188 7948 8192
rect 7884 8132 7888 8188
rect 7888 8132 7944 8188
rect 7944 8132 7948 8188
rect 7884 8128 7948 8132
rect 7964 8188 8028 8192
rect 7964 8132 7968 8188
rect 7968 8132 8024 8188
rect 8024 8132 8028 8188
rect 7964 8128 8028 8132
rect 8044 8188 8108 8192
rect 8044 8132 8048 8188
rect 8048 8132 8104 8188
rect 8104 8132 8108 8188
rect 8044 8128 8108 8132
rect 11506 8188 11570 8192
rect 11506 8132 11510 8188
rect 11510 8132 11566 8188
rect 11566 8132 11570 8188
rect 11506 8128 11570 8132
rect 11586 8188 11650 8192
rect 11586 8132 11590 8188
rect 11590 8132 11646 8188
rect 11646 8132 11650 8188
rect 11586 8128 11650 8132
rect 11666 8188 11730 8192
rect 11666 8132 11670 8188
rect 11670 8132 11726 8188
rect 11726 8132 11730 8188
rect 11666 8128 11730 8132
rect 11746 8188 11810 8192
rect 11746 8132 11750 8188
rect 11750 8132 11806 8188
rect 11806 8132 11810 8188
rect 11746 8128 11810 8132
rect 15208 8188 15272 8192
rect 15208 8132 15212 8188
rect 15212 8132 15268 8188
rect 15268 8132 15272 8188
rect 15208 8128 15272 8132
rect 15288 8188 15352 8192
rect 15288 8132 15292 8188
rect 15292 8132 15348 8188
rect 15348 8132 15352 8188
rect 15288 8128 15352 8132
rect 15368 8188 15432 8192
rect 15368 8132 15372 8188
rect 15372 8132 15428 8188
rect 15428 8132 15432 8188
rect 15368 8128 15432 8132
rect 15448 8188 15512 8192
rect 15448 8132 15452 8188
rect 15452 8132 15508 8188
rect 15508 8132 15512 8188
rect 15448 8128 15512 8132
rect 2251 7644 2315 7648
rect 2251 7588 2255 7644
rect 2255 7588 2311 7644
rect 2311 7588 2315 7644
rect 2251 7584 2315 7588
rect 2331 7644 2395 7648
rect 2331 7588 2335 7644
rect 2335 7588 2391 7644
rect 2391 7588 2395 7644
rect 2331 7584 2395 7588
rect 2411 7644 2475 7648
rect 2411 7588 2415 7644
rect 2415 7588 2471 7644
rect 2471 7588 2475 7644
rect 2411 7584 2475 7588
rect 2491 7644 2555 7648
rect 2491 7588 2495 7644
rect 2495 7588 2551 7644
rect 2551 7588 2555 7644
rect 2491 7584 2555 7588
rect 5953 7644 6017 7648
rect 5953 7588 5957 7644
rect 5957 7588 6013 7644
rect 6013 7588 6017 7644
rect 5953 7584 6017 7588
rect 6033 7644 6097 7648
rect 6033 7588 6037 7644
rect 6037 7588 6093 7644
rect 6093 7588 6097 7644
rect 6033 7584 6097 7588
rect 6113 7644 6177 7648
rect 6113 7588 6117 7644
rect 6117 7588 6173 7644
rect 6173 7588 6177 7644
rect 6113 7584 6177 7588
rect 6193 7644 6257 7648
rect 6193 7588 6197 7644
rect 6197 7588 6253 7644
rect 6253 7588 6257 7644
rect 6193 7584 6257 7588
rect 9655 7644 9719 7648
rect 9655 7588 9659 7644
rect 9659 7588 9715 7644
rect 9715 7588 9719 7644
rect 9655 7584 9719 7588
rect 9735 7644 9799 7648
rect 9735 7588 9739 7644
rect 9739 7588 9795 7644
rect 9795 7588 9799 7644
rect 9735 7584 9799 7588
rect 9815 7644 9879 7648
rect 9815 7588 9819 7644
rect 9819 7588 9875 7644
rect 9875 7588 9879 7644
rect 9815 7584 9879 7588
rect 9895 7644 9959 7648
rect 9895 7588 9899 7644
rect 9899 7588 9955 7644
rect 9955 7588 9959 7644
rect 9895 7584 9959 7588
rect 13357 7644 13421 7648
rect 13357 7588 13361 7644
rect 13361 7588 13417 7644
rect 13417 7588 13421 7644
rect 13357 7584 13421 7588
rect 13437 7644 13501 7648
rect 13437 7588 13441 7644
rect 13441 7588 13497 7644
rect 13497 7588 13501 7644
rect 13437 7584 13501 7588
rect 13517 7644 13581 7648
rect 13517 7588 13521 7644
rect 13521 7588 13577 7644
rect 13577 7588 13581 7644
rect 13517 7584 13581 7588
rect 13597 7644 13661 7648
rect 13597 7588 13601 7644
rect 13601 7588 13657 7644
rect 13657 7588 13661 7644
rect 13597 7584 13661 7588
rect 4102 7100 4166 7104
rect 4102 7044 4106 7100
rect 4106 7044 4162 7100
rect 4162 7044 4166 7100
rect 4102 7040 4166 7044
rect 4182 7100 4246 7104
rect 4182 7044 4186 7100
rect 4186 7044 4242 7100
rect 4242 7044 4246 7100
rect 4182 7040 4246 7044
rect 4262 7100 4326 7104
rect 4262 7044 4266 7100
rect 4266 7044 4322 7100
rect 4322 7044 4326 7100
rect 4262 7040 4326 7044
rect 4342 7100 4406 7104
rect 4342 7044 4346 7100
rect 4346 7044 4402 7100
rect 4402 7044 4406 7100
rect 4342 7040 4406 7044
rect 7804 7100 7868 7104
rect 7804 7044 7808 7100
rect 7808 7044 7864 7100
rect 7864 7044 7868 7100
rect 7804 7040 7868 7044
rect 7884 7100 7948 7104
rect 7884 7044 7888 7100
rect 7888 7044 7944 7100
rect 7944 7044 7948 7100
rect 7884 7040 7948 7044
rect 7964 7100 8028 7104
rect 7964 7044 7968 7100
rect 7968 7044 8024 7100
rect 8024 7044 8028 7100
rect 7964 7040 8028 7044
rect 8044 7100 8108 7104
rect 8044 7044 8048 7100
rect 8048 7044 8104 7100
rect 8104 7044 8108 7100
rect 8044 7040 8108 7044
rect 11506 7100 11570 7104
rect 11506 7044 11510 7100
rect 11510 7044 11566 7100
rect 11566 7044 11570 7100
rect 11506 7040 11570 7044
rect 11586 7100 11650 7104
rect 11586 7044 11590 7100
rect 11590 7044 11646 7100
rect 11646 7044 11650 7100
rect 11586 7040 11650 7044
rect 11666 7100 11730 7104
rect 11666 7044 11670 7100
rect 11670 7044 11726 7100
rect 11726 7044 11730 7100
rect 11666 7040 11730 7044
rect 11746 7100 11810 7104
rect 11746 7044 11750 7100
rect 11750 7044 11806 7100
rect 11806 7044 11810 7100
rect 11746 7040 11810 7044
rect 15208 7100 15272 7104
rect 15208 7044 15212 7100
rect 15212 7044 15268 7100
rect 15268 7044 15272 7100
rect 15208 7040 15272 7044
rect 15288 7100 15352 7104
rect 15288 7044 15292 7100
rect 15292 7044 15348 7100
rect 15348 7044 15352 7100
rect 15288 7040 15352 7044
rect 15368 7100 15432 7104
rect 15368 7044 15372 7100
rect 15372 7044 15428 7100
rect 15428 7044 15432 7100
rect 15368 7040 15432 7044
rect 15448 7100 15512 7104
rect 15448 7044 15452 7100
rect 15452 7044 15508 7100
rect 15508 7044 15512 7100
rect 15448 7040 15512 7044
rect 2251 6556 2315 6560
rect 2251 6500 2255 6556
rect 2255 6500 2311 6556
rect 2311 6500 2315 6556
rect 2251 6496 2315 6500
rect 2331 6556 2395 6560
rect 2331 6500 2335 6556
rect 2335 6500 2391 6556
rect 2391 6500 2395 6556
rect 2331 6496 2395 6500
rect 2411 6556 2475 6560
rect 2411 6500 2415 6556
rect 2415 6500 2471 6556
rect 2471 6500 2475 6556
rect 2411 6496 2475 6500
rect 2491 6556 2555 6560
rect 2491 6500 2495 6556
rect 2495 6500 2551 6556
rect 2551 6500 2555 6556
rect 2491 6496 2555 6500
rect 5953 6556 6017 6560
rect 5953 6500 5957 6556
rect 5957 6500 6013 6556
rect 6013 6500 6017 6556
rect 5953 6496 6017 6500
rect 6033 6556 6097 6560
rect 6033 6500 6037 6556
rect 6037 6500 6093 6556
rect 6093 6500 6097 6556
rect 6033 6496 6097 6500
rect 6113 6556 6177 6560
rect 6113 6500 6117 6556
rect 6117 6500 6173 6556
rect 6173 6500 6177 6556
rect 6113 6496 6177 6500
rect 6193 6556 6257 6560
rect 6193 6500 6197 6556
rect 6197 6500 6253 6556
rect 6253 6500 6257 6556
rect 6193 6496 6257 6500
rect 9655 6556 9719 6560
rect 9655 6500 9659 6556
rect 9659 6500 9715 6556
rect 9715 6500 9719 6556
rect 9655 6496 9719 6500
rect 9735 6556 9799 6560
rect 9735 6500 9739 6556
rect 9739 6500 9795 6556
rect 9795 6500 9799 6556
rect 9735 6496 9799 6500
rect 9815 6556 9879 6560
rect 9815 6500 9819 6556
rect 9819 6500 9875 6556
rect 9875 6500 9879 6556
rect 9815 6496 9879 6500
rect 9895 6556 9959 6560
rect 9895 6500 9899 6556
rect 9899 6500 9955 6556
rect 9955 6500 9959 6556
rect 9895 6496 9959 6500
rect 13357 6556 13421 6560
rect 13357 6500 13361 6556
rect 13361 6500 13417 6556
rect 13417 6500 13421 6556
rect 13357 6496 13421 6500
rect 13437 6556 13501 6560
rect 13437 6500 13441 6556
rect 13441 6500 13497 6556
rect 13497 6500 13501 6556
rect 13437 6496 13501 6500
rect 13517 6556 13581 6560
rect 13517 6500 13521 6556
rect 13521 6500 13577 6556
rect 13577 6500 13581 6556
rect 13517 6496 13581 6500
rect 13597 6556 13661 6560
rect 13597 6500 13601 6556
rect 13601 6500 13657 6556
rect 13657 6500 13661 6556
rect 13597 6496 13661 6500
rect 4102 6012 4166 6016
rect 4102 5956 4106 6012
rect 4106 5956 4162 6012
rect 4162 5956 4166 6012
rect 4102 5952 4166 5956
rect 4182 6012 4246 6016
rect 4182 5956 4186 6012
rect 4186 5956 4242 6012
rect 4242 5956 4246 6012
rect 4182 5952 4246 5956
rect 4262 6012 4326 6016
rect 4262 5956 4266 6012
rect 4266 5956 4322 6012
rect 4322 5956 4326 6012
rect 4262 5952 4326 5956
rect 4342 6012 4406 6016
rect 4342 5956 4346 6012
rect 4346 5956 4402 6012
rect 4402 5956 4406 6012
rect 4342 5952 4406 5956
rect 7804 6012 7868 6016
rect 7804 5956 7808 6012
rect 7808 5956 7864 6012
rect 7864 5956 7868 6012
rect 7804 5952 7868 5956
rect 7884 6012 7948 6016
rect 7884 5956 7888 6012
rect 7888 5956 7944 6012
rect 7944 5956 7948 6012
rect 7884 5952 7948 5956
rect 7964 6012 8028 6016
rect 7964 5956 7968 6012
rect 7968 5956 8024 6012
rect 8024 5956 8028 6012
rect 7964 5952 8028 5956
rect 8044 6012 8108 6016
rect 8044 5956 8048 6012
rect 8048 5956 8104 6012
rect 8104 5956 8108 6012
rect 8044 5952 8108 5956
rect 11506 6012 11570 6016
rect 11506 5956 11510 6012
rect 11510 5956 11566 6012
rect 11566 5956 11570 6012
rect 11506 5952 11570 5956
rect 11586 6012 11650 6016
rect 11586 5956 11590 6012
rect 11590 5956 11646 6012
rect 11646 5956 11650 6012
rect 11586 5952 11650 5956
rect 11666 6012 11730 6016
rect 11666 5956 11670 6012
rect 11670 5956 11726 6012
rect 11726 5956 11730 6012
rect 11666 5952 11730 5956
rect 11746 6012 11810 6016
rect 11746 5956 11750 6012
rect 11750 5956 11806 6012
rect 11806 5956 11810 6012
rect 11746 5952 11810 5956
rect 15208 6012 15272 6016
rect 15208 5956 15212 6012
rect 15212 5956 15268 6012
rect 15268 5956 15272 6012
rect 15208 5952 15272 5956
rect 15288 6012 15352 6016
rect 15288 5956 15292 6012
rect 15292 5956 15348 6012
rect 15348 5956 15352 6012
rect 15288 5952 15352 5956
rect 15368 6012 15432 6016
rect 15368 5956 15372 6012
rect 15372 5956 15428 6012
rect 15428 5956 15432 6012
rect 15368 5952 15432 5956
rect 15448 6012 15512 6016
rect 15448 5956 15452 6012
rect 15452 5956 15508 6012
rect 15508 5956 15512 6012
rect 15448 5952 15512 5956
rect 2251 5468 2315 5472
rect 2251 5412 2255 5468
rect 2255 5412 2311 5468
rect 2311 5412 2315 5468
rect 2251 5408 2315 5412
rect 2331 5468 2395 5472
rect 2331 5412 2335 5468
rect 2335 5412 2391 5468
rect 2391 5412 2395 5468
rect 2331 5408 2395 5412
rect 2411 5468 2475 5472
rect 2411 5412 2415 5468
rect 2415 5412 2471 5468
rect 2471 5412 2475 5468
rect 2411 5408 2475 5412
rect 2491 5468 2555 5472
rect 2491 5412 2495 5468
rect 2495 5412 2551 5468
rect 2551 5412 2555 5468
rect 2491 5408 2555 5412
rect 5953 5468 6017 5472
rect 5953 5412 5957 5468
rect 5957 5412 6013 5468
rect 6013 5412 6017 5468
rect 5953 5408 6017 5412
rect 6033 5468 6097 5472
rect 6033 5412 6037 5468
rect 6037 5412 6093 5468
rect 6093 5412 6097 5468
rect 6033 5408 6097 5412
rect 6113 5468 6177 5472
rect 6113 5412 6117 5468
rect 6117 5412 6173 5468
rect 6173 5412 6177 5468
rect 6113 5408 6177 5412
rect 6193 5468 6257 5472
rect 6193 5412 6197 5468
rect 6197 5412 6253 5468
rect 6253 5412 6257 5468
rect 6193 5408 6257 5412
rect 9655 5468 9719 5472
rect 9655 5412 9659 5468
rect 9659 5412 9715 5468
rect 9715 5412 9719 5468
rect 9655 5408 9719 5412
rect 9735 5468 9799 5472
rect 9735 5412 9739 5468
rect 9739 5412 9795 5468
rect 9795 5412 9799 5468
rect 9735 5408 9799 5412
rect 9815 5468 9879 5472
rect 9815 5412 9819 5468
rect 9819 5412 9875 5468
rect 9875 5412 9879 5468
rect 9815 5408 9879 5412
rect 9895 5468 9959 5472
rect 9895 5412 9899 5468
rect 9899 5412 9955 5468
rect 9955 5412 9959 5468
rect 9895 5408 9959 5412
rect 13357 5468 13421 5472
rect 13357 5412 13361 5468
rect 13361 5412 13417 5468
rect 13417 5412 13421 5468
rect 13357 5408 13421 5412
rect 13437 5468 13501 5472
rect 13437 5412 13441 5468
rect 13441 5412 13497 5468
rect 13497 5412 13501 5468
rect 13437 5408 13501 5412
rect 13517 5468 13581 5472
rect 13517 5412 13521 5468
rect 13521 5412 13577 5468
rect 13577 5412 13581 5468
rect 13517 5408 13581 5412
rect 13597 5468 13661 5472
rect 13597 5412 13601 5468
rect 13601 5412 13657 5468
rect 13657 5412 13661 5468
rect 13597 5408 13661 5412
rect 4102 4924 4166 4928
rect 4102 4868 4106 4924
rect 4106 4868 4162 4924
rect 4162 4868 4166 4924
rect 4102 4864 4166 4868
rect 4182 4924 4246 4928
rect 4182 4868 4186 4924
rect 4186 4868 4242 4924
rect 4242 4868 4246 4924
rect 4182 4864 4246 4868
rect 4262 4924 4326 4928
rect 4262 4868 4266 4924
rect 4266 4868 4322 4924
rect 4322 4868 4326 4924
rect 4262 4864 4326 4868
rect 4342 4924 4406 4928
rect 4342 4868 4346 4924
rect 4346 4868 4402 4924
rect 4402 4868 4406 4924
rect 4342 4864 4406 4868
rect 7804 4924 7868 4928
rect 7804 4868 7808 4924
rect 7808 4868 7864 4924
rect 7864 4868 7868 4924
rect 7804 4864 7868 4868
rect 7884 4924 7948 4928
rect 7884 4868 7888 4924
rect 7888 4868 7944 4924
rect 7944 4868 7948 4924
rect 7884 4864 7948 4868
rect 7964 4924 8028 4928
rect 7964 4868 7968 4924
rect 7968 4868 8024 4924
rect 8024 4868 8028 4924
rect 7964 4864 8028 4868
rect 8044 4924 8108 4928
rect 8044 4868 8048 4924
rect 8048 4868 8104 4924
rect 8104 4868 8108 4924
rect 8044 4864 8108 4868
rect 11506 4924 11570 4928
rect 11506 4868 11510 4924
rect 11510 4868 11566 4924
rect 11566 4868 11570 4924
rect 11506 4864 11570 4868
rect 11586 4924 11650 4928
rect 11586 4868 11590 4924
rect 11590 4868 11646 4924
rect 11646 4868 11650 4924
rect 11586 4864 11650 4868
rect 11666 4924 11730 4928
rect 11666 4868 11670 4924
rect 11670 4868 11726 4924
rect 11726 4868 11730 4924
rect 11666 4864 11730 4868
rect 11746 4924 11810 4928
rect 11746 4868 11750 4924
rect 11750 4868 11806 4924
rect 11806 4868 11810 4924
rect 11746 4864 11810 4868
rect 15208 4924 15272 4928
rect 15208 4868 15212 4924
rect 15212 4868 15268 4924
rect 15268 4868 15272 4924
rect 15208 4864 15272 4868
rect 15288 4924 15352 4928
rect 15288 4868 15292 4924
rect 15292 4868 15348 4924
rect 15348 4868 15352 4924
rect 15288 4864 15352 4868
rect 15368 4924 15432 4928
rect 15368 4868 15372 4924
rect 15372 4868 15428 4924
rect 15428 4868 15432 4924
rect 15368 4864 15432 4868
rect 15448 4924 15512 4928
rect 15448 4868 15452 4924
rect 15452 4868 15508 4924
rect 15508 4868 15512 4924
rect 15448 4864 15512 4868
rect 2251 4380 2315 4384
rect 2251 4324 2255 4380
rect 2255 4324 2311 4380
rect 2311 4324 2315 4380
rect 2251 4320 2315 4324
rect 2331 4380 2395 4384
rect 2331 4324 2335 4380
rect 2335 4324 2391 4380
rect 2391 4324 2395 4380
rect 2331 4320 2395 4324
rect 2411 4380 2475 4384
rect 2411 4324 2415 4380
rect 2415 4324 2471 4380
rect 2471 4324 2475 4380
rect 2411 4320 2475 4324
rect 2491 4380 2555 4384
rect 2491 4324 2495 4380
rect 2495 4324 2551 4380
rect 2551 4324 2555 4380
rect 2491 4320 2555 4324
rect 5953 4380 6017 4384
rect 5953 4324 5957 4380
rect 5957 4324 6013 4380
rect 6013 4324 6017 4380
rect 5953 4320 6017 4324
rect 6033 4380 6097 4384
rect 6033 4324 6037 4380
rect 6037 4324 6093 4380
rect 6093 4324 6097 4380
rect 6033 4320 6097 4324
rect 6113 4380 6177 4384
rect 6113 4324 6117 4380
rect 6117 4324 6173 4380
rect 6173 4324 6177 4380
rect 6113 4320 6177 4324
rect 6193 4380 6257 4384
rect 6193 4324 6197 4380
rect 6197 4324 6253 4380
rect 6253 4324 6257 4380
rect 6193 4320 6257 4324
rect 9655 4380 9719 4384
rect 9655 4324 9659 4380
rect 9659 4324 9715 4380
rect 9715 4324 9719 4380
rect 9655 4320 9719 4324
rect 9735 4380 9799 4384
rect 9735 4324 9739 4380
rect 9739 4324 9795 4380
rect 9795 4324 9799 4380
rect 9735 4320 9799 4324
rect 9815 4380 9879 4384
rect 9815 4324 9819 4380
rect 9819 4324 9875 4380
rect 9875 4324 9879 4380
rect 9815 4320 9879 4324
rect 9895 4380 9959 4384
rect 9895 4324 9899 4380
rect 9899 4324 9955 4380
rect 9955 4324 9959 4380
rect 9895 4320 9959 4324
rect 13357 4380 13421 4384
rect 13357 4324 13361 4380
rect 13361 4324 13417 4380
rect 13417 4324 13421 4380
rect 13357 4320 13421 4324
rect 13437 4380 13501 4384
rect 13437 4324 13441 4380
rect 13441 4324 13497 4380
rect 13497 4324 13501 4380
rect 13437 4320 13501 4324
rect 13517 4380 13581 4384
rect 13517 4324 13521 4380
rect 13521 4324 13577 4380
rect 13577 4324 13581 4380
rect 13517 4320 13581 4324
rect 13597 4380 13661 4384
rect 13597 4324 13601 4380
rect 13601 4324 13657 4380
rect 13657 4324 13661 4380
rect 13597 4320 13661 4324
rect 4102 3836 4166 3840
rect 4102 3780 4106 3836
rect 4106 3780 4162 3836
rect 4162 3780 4166 3836
rect 4102 3776 4166 3780
rect 4182 3836 4246 3840
rect 4182 3780 4186 3836
rect 4186 3780 4242 3836
rect 4242 3780 4246 3836
rect 4182 3776 4246 3780
rect 4262 3836 4326 3840
rect 4262 3780 4266 3836
rect 4266 3780 4322 3836
rect 4322 3780 4326 3836
rect 4262 3776 4326 3780
rect 4342 3836 4406 3840
rect 4342 3780 4346 3836
rect 4346 3780 4402 3836
rect 4402 3780 4406 3836
rect 4342 3776 4406 3780
rect 7804 3836 7868 3840
rect 7804 3780 7808 3836
rect 7808 3780 7864 3836
rect 7864 3780 7868 3836
rect 7804 3776 7868 3780
rect 7884 3836 7948 3840
rect 7884 3780 7888 3836
rect 7888 3780 7944 3836
rect 7944 3780 7948 3836
rect 7884 3776 7948 3780
rect 7964 3836 8028 3840
rect 7964 3780 7968 3836
rect 7968 3780 8024 3836
rect 8024 3780 8028 3836
rect 7964 3776 8028 3780
rect 8044 3836 8108 3840
rect 8044 3780 8048 3836
rect 8048 3780 8104 3836
rect 8104 3780 8108 3836
rect 8044 3776 8108 3780
rect 11506 3836 11570 3840
rect 11506 3780 11510 3836
rect 11510 3780 11566 3836
rect 11566 3780 11570 3836
rect 11506 3776 11570 3780
rect 11586 3836 11650 3840
rect 11586 3780 11590 3836
rect 11590 3780 11646 3836
rect 11646 3780 11650 3836
rect 11586 3776 11650 3780
rect 11666 3836 11730 3840
rect 11666 3780 11670 3836
rect 11670 3780 11726 3836
rect 11726 3780 11730 3836
rect 11666 3776 11730 3780
rect 11746 3836 11810 3840
rect 11746 3780 11750 3836
rect 11750 3780 11806 3836
rect 11806 3780 11810 3836
rect 11746 3776 11810 3780
rect 15208 3836 15272 3840
rect 15208 3780 15212 3836
rect 15212 3780 15268 3836
rect 15268 3780 15272 3836
rect 15208 3776 15272 3780
rect 15288 3836 15352 3840
rect 15288 3780 15292 3836
rect 15292 3780 15348 3836
rect 15348 3780 15352 3836
rect 15288 3776 15352 3780
rect 15368 3836 15432 3840
rect 15368 3780 15372 3836
rect 15372 3780 15428 3836
rect 15428 3780 15432 3836
rect 15368 3776 15432 3780
rect 15448 3836 15512 3840
rect 15448 3780 15452 3836
rect 15452 3780 15508 3836
rect 15508 3780 15512 3836
rect 15448 3776 15512 3780
rect 2251 3292 2315 3296
rect 2251 3236 2255 3292
rect 2255 3236 2311 3292
rect 2311 3236 2315 3292
rect 2251 3232 2315 3236
rect 2331 3292 2395 3296
rect 2331 3236 2335 3292
rect 2335 3236 2391 3292
rect 2391 3236 2395 3292
rect 2331 3232 2395 3236
rect 2411 3292 2475 3296
rect 2411 3236 2415 3292
rect 2415 3236 2471 3292
rect 2471 3236 2475 3292
rect 2411 3232 2475 3236
rect 2491 3292 2555 3296
rect 2491 3236 2495 3292
rect 2495 3236 2551 3292
rect 2551 3236 2555 3292
rect 2491 3232 2555 3236
rect 5953 3292 6017 3296
rect 5953 3236 5957 3292
rect 5957 3236 6013 3292
rect 6013 3236 6017 3292
rect 5953 3232 6017 3236
rect 6033 3292 6097 3296
rect 6033 3236 6037 3292
rect 6037 3236 6093 3292
rect 6093 3236 6097 3292
rect 6033 3232 6097 3236
rect 6113 3292 6177 3296
rect 6113 3236 6117 3292
rect 6117 3236 6173 3292
rect 6173 3236 6177 3292
rect 6113 3232 6177 3236
rect 6193 3292 6257 3296
rect 6193 3236 6197 3292
rect 6197 3236 6253 3292
rect 6253 3236 6257 3292
rect 6193 3232 6257 3236
rect 9655 3292 9719 3296
rect 9655 3236 9659 3292
rect 9659 3236 9715 3292
rect 9715 3236 9719 3292
rect 9655 3232 9719 3236
rect 9735 3292 9799 3296
rect 9735 3236 9739 3292
rect 9739 3236 9795 3292
rect 9795 3236 9799 3292
rect 9735 3232 9799 3236
rect 9815 3292 9879 3296
rect 9815 3236 9819 3292
rect 9819 3236 9875 3292
rect 9875 3236 9879 3292
rect 9815 3232 9879 3236
rect 9895 3292 9959 3296
rect 9895 3236 9899 3292
rect 9899 3236 9955 3292
rect 9955 3236 9959 3292
rect 9895 3232 9959 3236
rect 13357 3292 13421 3296
rect 13357 3236 13361 3292
rect 13361 3236 13417 3292
rect 13417 3236 13421 3292
rect 13357 3232 13421 3236
rect 13437 3292 13501 3296
rect 13437 3236 13441 3292
rect 13441 3236 13497 3292
rect 13497 3236 13501 3292
rect 13437 3232 13501 3236
rect 13517 3292 13581 3296
rect 13517 3236 13521 3292
rect 13521 3236 13577 3292
rect 13577 3236 13581 3292
rect 13517 3232 13581 3236
rect 13597 3292 13661 3296
rect 13597 3236 13601 3292
rect 13601 3236 13657 3292
rect 13657 3236 13661 3292
rect 13597 3232 13661 3236
rect 4102 2748 4166 2752
rect 4102 2692 4106 2748
rect 4106 2692 4162 2748
rect 4162 2692 4166 2748
rect 4102 2688 4166 2692
rect 4182 2748 4246 2752
rect 4182 2692 4186 2748
rect 4186 2692 4242 2748
rect 4242 2692 4246 2748
rect 4182 2688 4246 2692
rect 4262 2748 4326 2752
rect 4262 2692 4266 2748
rect 4266 2692 4322 2748
rect 4322 2692 4326 2748
rect 4262 2688 4326 2692
rect 4342 2748 4406 2752
rect 4342 2692 4346 2748
rect 4346 2692 4402 2748
rect 4402 2692 4406 2748
rect 4342 2688 4406 2692
rect 7804 2748 7868 2752
rect 7804 2692 7808 2748
rect 7808 2692 7864 2748
rect 7864 2692 7868 2748
rect 7804 2688 7868 2692
rect 7884 2748 7948 2752
rect 7884 2692 7888 2748
rect 7888 2692 7944 2748
rect 7944 2692 7948 2748
rect 7884 2688 7948 2692
rect 7964 2748 8028 2752
rect 7964 2692 7968 2748
rect 7968 2692 8024 2748
rect 8024 2692 8028 2748
rect 7964 2688 8028 2692
rect 8044 2748 8108 2752
rect 8044 2692 8048 2748
rect 8048 2692 8104 2748
rect 8104 2692 8108 2748
rect 8044 2688 8108 2692
rect 11506 2748 11570 2752
rect 11506 2692 11510 2748
rect 11510 2692 11566 2748
rect 11566 2692 11570 2748
rect 11506 2688 11570 2692
rect 11586 2748 11650 2752
rect 11586 2692 11590 2748
rect 11590 2692 11646 2748
rect 11646 2692 11650 2748
rect 11586 2688 11650 2692
rect 11666 2748 11730 2752
rect 11666 2692 11670 2748
rect 11670 2692 11726 2748
rect 11726 2692 11730 2748
rect 11666 2688 11730 2692
rect 11746 2748 11810 2752
rect 11746 2692 11750 2748
rect 11750 2692 11806 2748
rect 11806 2692 11810 2748
rect 11746 2688 11810 2692
rect 15208 2748 15272 2752
rect 15208 2692 15212 2748
rect 15212 2692 15268 2748
rect 15268 2692 15272 2748
rect 15208 2688 15272 2692
rect 15288 2748 15352 2752
rect 15288 2692 15292 2748
rect 15292 2692 15348 2748
rect 15348 2692 15352 2748
rect 15288 2688 15352 2692
rect 15368 2748 15432 2752
rect 15368 2692 15372 2748
rect 15372 2692 15428 2748
rect 15428 2692 15432 2748
rect 15368 2688 15432 2692
rect 15448 2748 15512 2752
rect 15448 2692 15452 2748
rect 15452 2692 15508 2748
rect 15508 2692 15512 2748
rect 15448 2688 15512 2692
rect 2251 2204 2315 2208
rect 2251 2148 2255 2204
rect 2255 2148 2311 2204
rect 2311 2148 2315 2204
rect 2251 2144 2315 2148
rect 2331 2204 2395 2208
rect 2331 2148 2335 2204
rect 2335 2148 2391 2204
rect 2391 2148 2395 2204
rect 2331 2144 2395 2148
rect 2411 2204 2475 2208
rect 2411 2148 2415 2204
rect 2415 2148 2471 2204
rect 2471 2148 2475 2204
rect 2411 2144 2475 2148
rect 2491 2204 2555 2208
rect 2491 2148 2495 2204
rect 2495 2148 2551 2204
rect 2551 2148 2555 2204
rect 2491 2144 2555 2148
rect 5953 2204 6017 2208
rect 5953 2148 5957 2204
rect 5957 2148 6013 2204
rect 6013 2148 6017 2204
rect 5953 2144 6017 2148
rect 6033 2204 6097 2208
rect 6033 2148 6037 2204
rect 6037 2148 6093 2204
rect 6093 2148 6097 2204
rect 6033 2144 6097 2148
rect 6113 2204 6177 2208
rect 6113 2148 6117 2204
rect 6117 2148 6173 2204
rect 6173 2148 6177 2204
rect 6113 2144 6177 2148
rect 6193 2204 6257 2208
rect 6193 2148 6197 2204
rect 6197 2148 6253 2204
rect 6253 2148 6257 2204
rect 6193 2144 6257 2148
rect 9655 2204 9719 2208
rect 9655 2148 9659 2204
rect 9659 2148 9715 2204
rect 9715 2148 9719 2204
rect 9655 2144 9719 2148
rect 9735 2204 9799 2208
rect 9735 2148 9739 2204
rect 9739 2148 9795 2204
rect 9795 2148 9799 2204
rect 9735 2144 9799 2148
rect 9815 2204 9879 2208
rect 9815 2148 9819 2204
rect 9819 2148 9875 2204
rect 9875 2148 9879 2204
rect 9815 2144 9879 2148
rect 9895 2204 9959 2208
rect 9895 2148 9899 2204
rect 9899 2148 9955 2204
rect 9955 2148 9959 2204
rect 9895 2144 9959 2148
rect 13357 2204 13421 2208
rect 13357 2148 13361 2204
rect 13361 2148 13417 2204
rect 13417 2148 13421 2204
rect 13357 2144 13421 2148
rect 13437 2204 13501 2208
rect 13437 2148 13441 2204
rect 13441 2148 13497 2204
rect 13497 2148 13501 2204
rect 13437 2144 13501 2148
rect 13517 2204 13581 2208
rect 13517 2148 13521 2204
rect 13521 2148 13577 2204
rect 13577 2148 13581 2204
rect 13517 2144 13581 2148
rect 13597 2204 13661 2208
rect 13597 2148 13601 2204
rect 13601 2148 13657 2204
rect 13657 2148 13661 2204
rect 13597 2144 13661 2148
rect 4102 1660 4166 1664
rect 4102 1604 4106 1660
rect 4106 1604 4162 1660
rect 4162 1604 4166 1660
rect 4102 1600 4166 1604
rect 4182 1660 4246 1664
rect 4182 1604 4186 1660
rect 4186 1604 4242 1660
rect 4242 1604 4246 1660
rect 4182 1600 4246 1604
rect 4262 1660 4326 1664
rect 4262 1604 4266 1660
rect 4266 1604 4322 1660
rect 4322 1604 4326 1660
rect 4262 1600 4326 1604
rect 4342 1660 4406 1664
rect 4342 1604 4346 1660
rect 4346 1604 4402 1660
rect 4402 1604 4406 1660
rect 4342 1600 4406 1604
rect 7804 1660 7868 1664
rect 7804 1604 7808 1660
rect 7808 1604 7864 1660
rect 7864 1604 7868 1660
rect 7804 1600 7868 1604
rect 7884 1660 7948 1664
rect 7884 1604 7888 1660
rect 7888 1604 7944 1660
rect 7944 1604 7948 1660
rect 7884 1600 7948 1604
rect 7964 1660 8028 1664
rect 7964 1604 7968 1660
rect 7968 1604 8024 1660
rect 8024 1604 8028 1660
rect 7964 1600 8028 1604
rect 8044 1660 8108 1664
rect 8044 1604 8048 1660
rect 8048 1604 8104 1660
rect 8104 1604 8108 1660
rect 8044 1600 8108 1604
rect 11506 1660 11570 1664
rect 11506 1604 11510 1660
rect 11510 1604 11566 1660
rect 11566 1604 11570 1660
rect 11506 1600 11570 1604
rect 11586 1660 11650 1664
rect 11586 1604 11590 1660
rect 11590 1604 11646 1660
rect 11646 1604 11650 1660
rect 11586 1600 11650 1604
rect 11666 1660 11730 1664
rect 11666 1604 11670 1660
rect 11670 1604 11726 1660
rect 11726 1604 11730 1660
rect 11666 1600 11730 1604
rect 11746 1660 11810 1664
rect 11746 1604 11750 1660
rect 11750 1604 11806 1660
rect 11806 1604 11810 1660
rect 11746 1600 11810 1604
rect 15208 1660 15272 1664
rect 15208 1604 15212 1660
rect 15212 1604 15268 1660
rect 15268 1604 15272 1660
rect 15208 1600 15272 1604
rect 15288 1660 15352 1664
rect 15288 1604 15292 1660
rect 15292 1604 15348 1660
rect 15348 1604 15352 1660
rect 15288 1600 15352 1604
rect 15368 1660 15432 1664
rect 15368 1604 15372 1660
rect 15372 1604 15428 1660
rect 15428 1604 15432 1660
rect 15368 1600 15432 1604
rect 15448 1660 15512 1664
rect 15448 1604 15452 1660
rect 15452 1604 15508 1660
rect 15508 1604 15512 1660
rect 15448 1600 15512 1604
rect 2251 1116 2315 1120
rect 2251 1060 2255 1116
rect 2255 1060 2311 1116
rect 2311 1060 2315 1116
rect 2251 1056 2315 1060
rect 2331 1116 2395 1120
rect 2331 1060 2335 1116
rect 2335 1060 2391 1116
rect 2391 1060 2395 1116
rect 2331 1056 2395 1060
rect 2411 1116 2475 1120
rect 2411 1060 2415 1116
rect 2415 1060 2471 1116
rect 2471 1060 2475 1116
rect 2411 1056 2475 1060
rect 2491 1116 2555 1120
rect 2491 1060 2495 1116
rect 2495 1060 2551 1116
rect 2551 1060 2555 1116
rect 2491 1056 2555 1060
rect 5953 1116 6017 1120
rect 5953 1060 5957 1116
rect 5957 1060 6013 1116
rect 6013 1060 6017 1116
rect 5953 1056 6017 1060
rect 6033 1116 6097 1120
rect 6033 1060 6037 1116
rect 6037 1060 6093 1116
rect 6093 1060 6097 1116
rect 6033 1056 6097 1060
rect 6113 1116 6177 1120
rect 6113 1060 6117 1116
rect 6117 1060 6173 1116
rect 6173 1060 6177 1116
rect 6113 1056 6177 1060
rect 6193 1116 6257 1120
rect 6193 1060 6197 1116
rect 6197 1060 6253 1116
rect 6253 1060 6257 1116
rect 6193 1056 6257 1060
rect 9655 1116 9719 1120
rect 9655 1060 9659 1116
rect 9659 1060 9715 1116
rect 9715 1060 9719 1116
rect 9655 1056 9719 1060
rect 9735 1116 9799 1120
rect 9735 1060 9739 1116
rect 9739 1060 9795 1116
rect 9795 1060 9799 1116
rect 9735 1056 9799 1060
rect 9815 1116 9879 1120
rect 9815 1060 9819 1116
rect 9819 1060 9875 1116
rect 9875 1060 9879 1116
rect 9815 1056 9879 1060
rect 9895 1116 9959 1120
rect 9895 1060 9899 1116
rect 9899 1060 9955 1116
rect 9955 1060 9959 1116
rect 9895 1056 9959 1060
rect 13357 1116 13421 1120
rect 13357 1060 13361 1116
rect 13361 1060 13417 1116
rect 13417 1060 13421 1116
rect 13357 1056 13421 1060
rect 13437 1116 13501 1120
rect 13437 1060 13441 1116
rect 13441 1060 13497 1116
rect 13497 1060 13501 1116
rect 13437 1056 13501 1060
rect 13517 1116 13581 1120
rect 13517 1060 13521 1116
rect 13521 1060 13577 1116
rect 13577 1060 13581 1116
rect 13517 1056 13581 1060
rect 13597 1116 13661 1120
rect 13597 1060 13601 1116
rect 13601 1060 13657 1116
rect 13657 1060 13661 1116
rect 13597 1056 13661 1060
rect 4102 572 4166 576
rect 4102 516 4106 572
rect 4106 516 4162 572
rect 4162 516 4166 572
rect 4102 512 4166 516
rect 4182 572 4246 576
rect 4182 516 4186 572
rect 4186 516 4242 572
rect 4242 516 4246 572
rect 4182 512 4246 516
rect 4262 572 4326 576
rect 4262 516 4266 572
rect 4266 516 4322 572
rect 4322 516 4326 572
rect 4262 512 4326 516
rect 4342 572 4406 576
rect 4342 516 4346 572
rect 4346 516 4402 572
rect 4402 516 4406 572
rect 4342 512 4406 516
rect 7804 572 7868 576
rect 7804 516 7808 572
rect 7808 516 7864 572
rect 7864 516 7868 572
rect 7804 512 7868 516
rect 7884 572 7948 576
rect 7884 516 7888 572
rect 7888 516 7944 572
rect 7944 516 7948 572
rect 7884 512 7948 516
rect 7964 572 8028 576
rect 7964 516 7968 572
rect 7968 516 8024 572
rect 8024 516 8028 572
rect 7964 512 8028 516
rect 8044 572 8108 576
rect 8044 516 8048 572
rect 8048 516 8104 572
rect 8104 516 8108 572
rect 8044 512 8108 516
rect 11506 572 11570 576
rect 11506 516 11510 572
rect 11510 516 11566 572
rect 11566 516 11570 572
rect 11506 512 11570 516
rect 11586 572 11650 576
rect 11586 516 11590 572
rect 11590 516 11646 572
rect 11646 516 11650 572
rect 11586 512 11650 516
rect 11666 572 11730 576
rect 11666 516 11670 572
rect 11670 516 11726 572
rect 11726 516 11730 572
rect 11666 512 11730 516
rect 11746 572 11810 576
rect 11746 516 11750 572
rect 11750 516 11806 572
rect 11806 516 11810 572
rect 11746 512 11810 516
rect 15208 572 15272 576
rect 15208 516 15212 572
rect 15212 516 15268 572
rect 15268 516 15272 572
rect 15208 512 15272 516
rect 15288 572 15352 576
rect 15288 516 15292 572
rect 15292 516 15348 572
rect 15348 516 15352 572
rect 15288 512 15352 516
rect 15368 572 15432 576
rect 15368 516 15372 572
rect 15372 516 15428 572
rect 15428 516 15432 572
rect 15368 512 15432 516
rect 15448 572 15512 576
rect 15448 516 15452 572
rect 15452 516 15508 572
rect 15508 516 15512 572
rect 15448 512 15512 516
<< metal4 >>
rect 2243 15264 2563 15280
rect 2243 15200 2251 15264
rect 2315 15200 2331 15264
rect 2395 15200 2411 15264
rect 2475 15200 2491 15264
rect 2555 15200 2563 15264
rect 2243 14176 2563 15200
rect 2243 14112 2251 14176
rect 2315 14112 2331 14176
rect 2395 14112 2411 14176
rect 2475 14112 2491 14176
rect 2555 14112 2563 14176
rect 2243 13088 2563 14112
rect 2243 13024 2251 13088
rect 2315 13024 2331 13088
rect 2395 13024 2411 13088
rect 2475 13024 2491 13088
rect 2555 13024 2563 13088
rect 2243 12000 2563 13024
rect 2243 11936 2251 12000
rect 2315 11936 2331 12000
rect 2395 11936 2411 12000
rect 2475 11936 2491 12000
rect 2555 11936 2563 12000
rect 2243 10912 2563 11936
rect 2243 10848 2251 10912
rect 2315 10848 2331 10912
rect 2395 10848 2411 10912
rect 2475 10848 2491 10912
rect 2555 10848 2563 10912
rect 2243 9824 2563 10848
rect 2243 9760 2251 9824
rect 2315 9760 2331 9824
rect 2395 9760 2411 9824
rect 2475 9760 2491 9824
rect 2555 9760 2563 9824
rect 2243 8736 2563 9760
rect 2243 8672 2251 8736
rect 2315 8672 2331 8736
rect 2395 8672 2411 8736
rect 2475 8672 2491 8736
rect 2555 8672 2563 8736
rect 2243 7648 2563 8672
rect 2243 7584 2251 7648
rect 2315 7584 2331 7648
rect 2395 7584 2411 7648
rect 2475 7584 2491 7648
rect 2555 7584 2563 7648
rect 2243 6560 2563 7584
rect 2243 6496 2251 6560
rect 2315 6496 2331 6560
rect 2395 6496 2411 6560
rect 2475 6496 2491 6560
rect 2555 6496 2563 6560
rect 2243 5472 2563 6496
rect 2243 5408 2251 5472
rect 2315 5408 2331 5472
rect 2395 5408 2411 5472
rect 2475 5408 2491 5472
rect 2555 5408 2563 5472
rect 2243 4384 2563 5408
rect 2243 4320 2251 4384
rect 2315 4320 2331 4384
rect 2395 4320 2411 4384
rect 2475 4320 2491 4384
rect 2555 4320 2563 4384
rect 2243 3296 2563 4320
rect 2243 3232 2251 3296
rect 2315 3232 2331 3296
rect 2395 3232 2411 3296
rect 2475 3232 2491 3296
rect 2555 3232 2563 3296
rect 2243 2208 2563 3232
rect 2243 2144 2251 2208
rect 2315 2144 2331 2208
rect 2395 2144 2411 2208
rect 2475 2144 2491 2208
rect 2555 2144 2563 2208
rect 2243 1120 2563 2144
rect 2243 1056 2251 1120
rect 2315 1056 2331 1120
rect 2395 1056 2411 1120
rect 2475 1056 2491 1120
rect 2555 1056 2563 1120
rect 2243 496 2563 1056
rect 4094 14720 4414 15280
rect 4094 14656 4102 14720
rect 4166 14656 4182 14720
rect 4246 14656 4262 14720
rect 4326 14656 4342 14720
rect 4406 14656 4414 14720
rect 4094 13632 4414 14656
rect 4094 13568 4102 13632
rect 4166 13568 4182 13632
rect 4246 13568 4262 13632
rect 4326 13568 4342 13632
rect 4406 13568 4414 13632
rect 4094 12544 4414 13568
rect 4094 12480 4102 12544
rect 4166 12480 4182 12544
rect 4246 12480 4262 12544
rect 4326 12480 4342 12544
rect 4406 12480 4414 12544
rect 4094 11456 4414 12480
rect 4094 11392 4102 11456
rect 4166 11392 4182 11456
rect 4246 11392 4262 11456
rect 4326 11392 4342 11456
rect 4406 11392 4414 11456
rect 4094 10368 4414 11392
rect 4094 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4342 10368
rect 4406 10304 4414 10368
rect 4094 9280 4414 10304
rect 4094 9216 4102 9280
rect 4166 9216 4182 9280
rect 4246 9216 4262 9280
rect 4326 9216 4342 9280
rect 4406 9216 4414 9280
rect 4094 8192 4414 9216
rect 4094 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4342 8192
rect 4406 8128 4414 8192
rect 4094 7104 4414 8128
rect 4094 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4342 7104
rect 4406 7040 4414 7104
rect 4094 6016 4414 7040
rect 4094 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4342 6016
rect 4406 5952 4414 6016
rect 4094 4928 4414 5952
rect 4094 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4342 4928
rect 4406 4864 4414 4928
rect 4094 3840 4414 4864
rect 4094 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4342 3840
rect 4406 3776 4414 3840
rect 4094 2752 4414 3776
rect 4094 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4342 2752
rect 4406 2688 4414 2752
rect 4094 1664 4414 2688
rect 4094 1600 4102 1664
rect 4166 1600 4182 1664
rect 4246 1600 4262 1664
rect 4326 1600 4342 1664
rect 4406 1600 4414 1664
rect 4094 576 4414 1600
rect 4094 512 4102 576
rect 4166 512 4182 576
rect 4246 512 4262 576
rect 4326 512 4342 576
rect 4406 512 4414 576
rect 4094 496 4414 512
rect 5945 15264 6265 15280
rect 5945 15200 5953 15264
rect 6017 15200 6033 15264
rect 6097 15200 6113 15264
rect 6177 15200 6193 15264
rect 6257 15200 6265 15264
rect 5945 14176 6265 15200
rect 5945 14112 5953 14176
rect 6017 14112 6033 14176
rect 6097 14112 6113 14176
rect 6177 14112 6193 14176
rect 6257 14112 6265 14176
rect 5945 13088 6265 14112
rect 5945 13024 5953 13088
rect 6017 13024 6033 13088
rect 6097 13024 6113 13088
rect 6177 13024 6193 13088
rect 6257 13024 6265 13088
rect 5945 12000 6265 13024
rect 5945 11936 5953 12000
rect 6017 11936 6033 12000
rect 6097 11936 6113 12000
rect 6177 11936 6193 12000
rect 6257 11936 6265 12000
rect 5945 10912 6265 11936
rect 5945 10848 5953 10912
rect 6017 10848 6033 10912
rect 6097 10848 6113 10912
rect 6177 10848 6193 10912
rect 6257 10848 6265 10912
rect 5945 9824 6265 10848
rect 5945 9760 5953 9824
rect 6017 9760 6033 9824
rect 6097 9760 6113 9824
rect 6177 9760 6193 9824
rect 6257 9760 6265 9824
rect 5945 8736 6265 9760
rect 5945 8672 5953 8736
rect 6017 8672 6033 8736
rect 6097 8672 6113 8736
rect 6177 8672 6193 8736
rect 6257 8672 6265 8736
rect 5945 7648 6265 8672
rect 5945 7584 5953 7648
rect 6017 7584 6033 7648
rect 6097 7584 6113 7648
rect 6177 7584 6193 7648
rect 6257 7584 6265 7648
rect 5945 6560 6265 7584
rect 5945 6496 5953 6560
rect 6017 6496 6033 6560
rect 6097 6496 6113 6560
rect 6177 6496 6193 6560
rect 6257 6496 6265 6560
rect 5945 5472 6265 6496
rect 5945 5408 5953 5472
rect 6017 5408 6033 5472
rect 6097 5408 6113 5472
rect 6177 5408 6193 5472
rect 6257 5408 6265 5472
rect 5945 4384 6265 5408
rect 5945 4320 5953 4384
rect 6017 4320 6033 4384
rect 6097 4320 6113 4384
rect 6177 4320 6193 4384
rect 6257 4320 6265 4384
rect 5945 3296 6265 4320
rect 5945 3232 5953 3296
rect 6017 3232 6033 3296
rect 6097 3232 6113 3296
rect 6177 3232 6193 3296
rect 6257 3232 6265 3296
rect 5945 2208 6265 3232
rect 5945 2144 5953 2208
rect 6017 2144 6033 2208
rect 6097 2144 6113 2208
rect 6177 2144 6193 2208
rect 6257 2144 6265 2208
rect 5945 1120 6265 2144
rect 5945 1056 5953 1120
rect 6017 1056 6033 1120
rect 6097 1056 6113 1120
rect 6177 1056 6193 1120
rect 6257 1056 6265 1120
rect 5945 496 6265 1056
rect 7796 14720 8116 15280
rect 7796 14656 7804 14720
rect 7868 14656 7884 14720
rect 7948 14656 7964 14720
rect 8028 14656 8044 14720
rect 8108 14656 8116 14720
rect 7796 13632 8116 14656
rect 7796 13568 7804 13632
rect 7868 13568 7884 13632
rect 7948 13568 7964 13632
rect 8028 13568 8044 13632
rect 8108 13568 8116 13632
rect 7796 12544 8116 13568
rect 7796 12480 7804 12544
rect 7868 12480 7884 12544
rect 7948 12480 7964 12544
rect 8028 12480 8044 12544
rect 8108 12480 8116 12544
rect 7796 11456 8116 12480
rect 7796 11392 7804 11456
rect 7868 11392 7884 11456
rect 7948 11392 7964 11456
rect 8028 11392 8044 11456
rect 8108 11392 8116 11456
rect 7796 10368 8116 11392
rect 7796 10304 7804 10368
rect 7868 10304 7884 10368
rect 7948 10304 7964 10368
rect 8028 10304 8044 10368
rect 8108 10304 8116 10368
rect 7796 9280 8116 10304
rect 7796 9216 7804 9280
rect 7868 9216 7884 9280
rect 7948 9216 7964 9280
rect 8028 9216 8044 9280
rect 8108 9216 8116 9280
rect 7796 8192 8116 9216
rect 7796 8128 7804 8192
rect 7868 8128 7884 8192
rect 7948 8128 7964 8192
rect 8028 8128 8044 8192
rect 8108 8128 8116 8192
rect 7796 7104 8116 8128
rect 7796 7040 7804 7104
rect 7868 7040 7884 7104
rect 7948 7040 7964 7104
rect 8028 7040 8044 7104
rect 8108 7040 8116 7104
rect 7796 6016 8116 7040
rect 7796 5952 7804 6016
rect 7868 5952 7884 6016
rect 7948 5952 7964 6016
rect 8028 5952 8044 6016
rect 8108 5952 8116 6016
rect 7796 4928 8116 5952
rect 7796 4864 7804 4928
rect 7868 4864 7884 4928
rect 7948 4864 7964 4928
rect 8028 4864 8044 4928
rect 8108 4864 8116 4928
rect 7796 3840 8116 4864
rect 7796 3776 7804 3840
rect 7868 3776 7884 3840
rect 7948 3776 7964 3840
rect 8028 3776 8044 3840
rect 8108 3776 8116 3840
rect 7796 2752 8116 3776
rect 7796 2688 7804 2752
rect 7868 2688 7884 2752
rect 7948 2688 7964 2752
rect 8028 2688 8044 2752
rect 8108 2688 8116 2752
rect 7796 1664 8116 2688
rect 7796 1600 7804 1664
rect 7868 1600 7884 1664
rect 7948 1600 7964 1664
rect 8028 1600 8044 1664
rect 8108 1600 8116 1664
rect 7796 576 8116 1600
rect 7796 512 7804 576
rect 7868 512 7884 576
rect 7948 512 7964 576
rect 8028 512 8044 576
rect 8108 512 8116 576
rect 7796 496 8116 512
rect 9647 15264 9967 15280
rect 9647 15200 9655 15264
rect 9719 15200 9735 15264
rect 9799 15200 9815 15264
rect 9879 15200 9895 15264
rect 9959 15200 9967 15264
rect 9647 14176 9967 15200
rect 9647 14112 9655 14176
rect 9719 14112 9735 14176
rect 9799 14112 9815 14176
rect 9879 14112 9895 14176
rect 9959 14112 9967 14176
rect 9647 13088 9967 14112
rect 9647 13024 9655 13088
rect 9719 13024 9735 13088
rect 9799 13024 9815 13088
rect 9879 13024 9895 13088
rect 9959 13024 9967 13088
rect 9647 12000 9967 13024
rect 9647 11936 9655 12000
rect 9719 11936 9735 12000
rect 9799 11936 9815 12000
rect 9879 11936 9895 12000
rect 9959 11936 9967 12000
rect 9647 10912 9967 11936
rect 9647 10848 9655 10912
rect 9719 10848 9735 10912
rect 9799 10848 9815 10912
rect 9879 10848 9895 10912
rect 9959 10848 9967 10912
rect 9647 9824 9967 10848
rect 9647 9760 9655 9824
rect 9719 9760 9735 9824
rect 9799 9760 9815 9824
rect 9879 9760 9895 9824
rect 9959 9760 9967 9824
rect 9647 8736 9967 9760
rect 9647 8672 9655 8736
rect 9719 8672 9735 8736
rect 9799 8672 9815 8736
rect 9879 8672 9895 8736
rect 9959 8672 9967 8736
rect 9647 7648 9967 8672
rect 9647 7584 9655 7648
rect 9719 7584 9735 7648
rect 9799 7584 9815 7648
rect 9879 7584 9895 7648
rect 9959 7584 9967 7648
rect 9647 6560 9967 7584
rect 9647 6496 9655 6560
rect 9719 6496 9735 6560
rect 9799 6496 9815 6560
rect 9879 6496 9895 6560
rect 9959 6496 9967 6560
rect 9647 5472 9967 6496
rect 9647 5408 9655 5472
rect 9719 5408 9735 5472
rect 9799 5408 9815 5472
rect 9879 5408 9895 5472
rect 9959 5408 9967 5472
rect 9647 4384 9967 5408
rect 9647 4320 9655 4384
rect 9719 4320 9735 4384
rect 9799 4320 9815 4384
rect 9879 4320 9895 4384
rect 9959 4320 9967 4384
rect 9647 3296 9967 4320
rect 9647 3232 9655 3296
rect 9719 3232 9735 3296
rect 9799 3232 9815 3296
rect 9879 3232 9895 3296
rect 9959 3232 9967 3296
rect 9647 2208 9967 3232
rect 9647 2144 9655 2208
rect 9719 2144 9735 2208
rect 9799 2144 9815 2208
rect 9879 2144 9895 2208
rect 9959 2144 9967 2208
rect 9647 1120 9967 2144
rect 9647 1056 9655 1120
rect 9719 1056 9735 1120
rect 9799 1056 9815 1120
rect 9879 1056 9895 1120
rect 9959 1056 9967 1120
rect 9647 496 9967 1056
rect 11498 14720 11818 15280
rect 11498 14656 11506 14720
rect 11570 14656 11586 14720
rect 11650 14656 11666 14720
rect 11730 14656 11746 14720
rect 11810 14656 11818 14720
rect 11498 13632 11818 14656
rect 11498 13568 11506 13632
rect 11570 13568 11586 13632
rect 11650 13568 11666 13632
rect 11730 13568 11746 13632
rect 11810 13568 11818 13632
rect 11498 12544 11818 13568
rect 11498 12480 11506 12544
rect 11570 12480 11586 12544
rect 11650 12480 11666 12544
rect 11730 12480 11746 12544
rect 11810 12480 11818 12544
rect 11498 11456 11818 12480
rect 11498 11392 11506 11456
rect 11570 11392 11586 11456
rect 11650 11392 11666 11456
rect 11730 11392 11746 11456
rect 11810 11392 11818 11456
rect 11498 10368 11818 11392
rect 11498 10304 11506 10368
rect 11570 10304 11586 10368
rect 11650 10304 11666 10368
rect 11730 10304 11746 10368
rect 11810 10304 11818 10368
rect 11498 9280 11818 10304
rect 11498 9216 11506 9280
rect 11570 9216 11586 9280
rect 11650 9216 11666 9280
rect 11730 9216 11746 9280
rect 11810 9216 11818 9280
rect 11498 8192 11818 9216
rect 11498 8128 11506 8192
rect 11570 8128 11586 8192
rect 11650 8128 11666 8192
rect 11730 8128 11746 8192
rect 11810 8128 11818 8192
rect 11498 7104 11818 8128
rect 11498 7040 11506 7104
rect 11570 7040 11586 7104
rect 11650 7040 11666 7104
rect 11730 7040 11746 7104
rect 11810 7040 11818 7104
rect 11498 6016 11818 7040
rect 11498 5952 11506 6016
rect 11570 5952 11586 6016
rect 11650 5952 11666 6016
rect 11730 5952 11746 6016
rect 11810 5952 11818 6016
rect 11498 4928 11818 5952
rect 11498 4864 11506 4928
rect 11570 4864 11586 4928
rect 11650 4864 11666 4928
rect 11730 4864 11746 4928
rect 11810 4864 11818 4928
rect 11498 3840 11818 4864
rect 11498 3776 11506 3840
rect 11570 3776 11586 3840
rect 11650 3776 11666 3840
rect 11730 3776 11746 3840
rect 11810 3776 11818 3840
rect 11498 2752 11818 3776
rect 11498 2688 11506 2752
rect 11570 2688 11586 2752
rect 11650 2688 11666 2752
rect 11730 2688 11746 2752
rect 11810 2688 11818 2752
rect 11498 1664 11818 2688
rect 11498 1600 11506 1664
rect 11570 1600 11586 1664
rect 11650 1600 11666 1664
rect 11730 1600 11746 1664
rect 11810 1600 11818 1664
rect 11498 576 11818 1600
rect 11498 512 11506 576
rect 11570 512 11586 576
rect 11650 512 11666 576
rect 11730 512 11746 576
rect 11810 512 11818 576
rect 11498 496 11818 512
rect 13349 15264 13669 15280
rect 13349 15200 13357 15264
rect 13421 15200 13437 15264
rect 13501 15200 13517 15264
rect 13581 15200 13597 15264
rect 13661 15200 13669 15264
rect 13349 14176 13669 15200
rect 13349 14112 13357 14176
rect 13421 14112 13437 14176
rect 13501 14112 13517 14176
rect 13581 14112 13597 14176
rect 13661 14112 13669 14176
rect 13349 13088 13669 14112
rect 13349 13024 13357 13088
rect 13421 13024 13437 13088
rect 13501 13024 13517 13088
rect 13581 13024 13597 13088
rect 13661 13024 13669 13088
rect 13349 12000 13669 13024
rect 13349 11936 13357 12000
rect 13421 11936 13437 12000
rect 13501 11936 13517 12000
rect 13581 11936 13597 12000
rect 13661 11936 13669 12000
rect 13349 10912 13669 11936
rect 13349 10848 13357 10912
rect 13421 10848 13437 10912
rect 13501 10848 13517 10912
rect 13581 10848 13597 10912
rect 13661 10848 13669 10912
rect 13349 9824 13669 10848
rect 13349 9760 13357 9824
rect 13421 9760 13437 9824
rect 13501 9760 13517 9824
rect 13581 9760 13597 9824
rect 13661 9760 13669 9824
rect 13349 8736 13669 9760
rect 13349 8672 13357 8736
rect 13421 8672 13437 8736
rect 13501 8672 13517 8736
rect 13581 8672 13597 8736
rect 13661 8672 13669 8736
rect 13349 7648 13669 8672
rect 13349 7584 13357 7648
rect 13421 7584 13437 7648
rect 13501 7584 13517 7648
rect 13581 7584 13597 7648
rect 13661 7584 13669 7648
rect 13349 6560 13669 7584
rect 13349 6496 13357 6560
rect 13421 6496 13437 6560
rect 13501 6496 13517 6560
rect 13581 6496 13597 6560
rect 13661 6496 13669 6560
rect 13349 5472 13669 6496
rect 13349 5408 13357 5472
rect 13421 5408 13437 5472
rect 13501 5408 13517 5472
rect 13581 5408 13597 5472
rect 13661 5408 13669 5472
rect 13349 4384 13669 5408
rect 13349 4320 13357 4384
rect 13421 4320 13437 4384
rect 13501 4320 13517 4384
rect 13581 4320 13597 4384
rect 13661 4320 13669 4384
rect 13349 3296 13669 4320
rect 13349 3232 13357 3296
rect 13421 3232 13437 3296
rect 13501 3232 13517 3296
rect 13581 3232 13597 3296
rect 13661 3232 13669 3296
rect 13349 2208 13669 3232
rect 13349 2144 13357 2208
rect 13421 2144 13437 2208
rect 13501 2144 13517 2208
rect 13581 2144 13597 2208
rect 13661 2144 13669 2208
rect 13349 1120 13669 2144
rect 13349 1056 13357 1120
rect 13421 1056 13437 1120
rect 13501 1056 13517 1120
rect 13581 1056 13597 1120
rect 13661 1056 13669 1120
rect 13349 496 13669 1056
rect 15200 14720 15520 15280
rect 15200 14656 15208 14720
rect 15272 14656 15288 14720
rect 15352 14656 15368 14720
rect 15432 14656 15448 14720
rect 15512 14656 15520 14720
rect 15200 13632 15520 14656
rect 15200 13568 15208 13632
rect 15272 13568 15288 13632
rect 15352 13568 15368 13632
rect 15432 13568 15448 13632
rect 15512 13568 15520 13632
rect 15200 12544 15520 13568
rect 15200 12480 15208 12544
rect 15272 12480 15288 12544
rect 15352 12480 15368 12544
rect 15432 12480 15448 12544
rect 15512 12480 15520 12544
rect 15200 11456 15520 12480
rect 15200 11392 15208 11456
rect 15272 11392 15288 11456
rect 15352 11392 15368 11456
rect 15432 11392 15448 11456
rect 15512 11392 15520 11456
rect 15200 10368 15520 11392
rect 15200 10304 15208 10368
rect 15272 10304 15288 10368
rect 15352 10304 15368 10368
rect 15432 10304 15448 10368
rect 15512 10304 15520 10368
rect 15200 9280 15520 10304
rect 15200 9216 15208 9280
rect 15272 9216 15288 9280
rect 15352 9216 15368 9280
rect 15432 9216 15448 9280
rect 15512 9216 15520 9280
rect 15200 8192 15520 9216
rect 15200 8128 15208 8192
rect 15272 8128 15288 8192
rect 15352 8128 15368 8192
rect 15432 8128 15448 8192
rect 15512 8128 15520 8192
rect 15200 7104 15520 8128
rect 15200 7040 15208 7104
rect 15272 7040 15288 7104
rect 15352 7040 15368 7104
rect 15432 7040 15448 7104
rect 15512 7040 15520 7104
rect 15200 6016 15520 7040
rect 15200 5952 15208 6016
rect 15272 5952 15288 6016
rect 15352 5952 15368 6016
rect 15432 5952 15448 6016
rect 15512 5952 15520 6016
rect 15200 4928 15520 5952
rect 15200 4864 15208 4928
rect 15272 4864 15288 4928
rect 15352 4864 15368 4928
rect 15432 4864 15448 4928
rect 15512 4864 15520 4928
rect 15200 3840 15520 4864
rect 15200 3776 15208 3840
rect 15272 3776 15288 3840
rect 15352 3776 15368 3840
rect 15432 3776 15448 3840
rect 15512 3776 15520 3840
rect 15200 2752 15520 3776
rect 15200 2688 15208 2752
rect 15272 2688 15288 2752
rect 15352 2688 15368 2752
rect 15432 2688 15448 2752
rect 15512 2688 15520 2752
rect 15200 1664 15520 2688
rect 15200 1600 15208 1664
rect 15272 1600 15288 1664
rect 15352 1600 15368 1664
rect 15432 1600 15448 1664
rect 15512 1600 15520 1664
rect 15200 576 15520 1600
rect 15200 512 15208 576
rect 15272 512 15288 576
rect 15352 512 15368 576
rect 15432 512 15448 576
rect 15512 512 15520 576
rect 15200 496 15520 512
use sky130_fd_sc_hd__mux2_1  _30_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10028 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _31_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14536 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _32_
timestamp 1688980957
transform 1 0 11868 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _33_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11500 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _34_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4876 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _35_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _36_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _37_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6164 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _38_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5060 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _39_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8832 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _40_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9476 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _41_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6256 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _42_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7728 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _43_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6624 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _44_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7912 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _45_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6900 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _46_
timestamp 1688980957
transform -1 0 10304 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _47_
timestamp 1688980957
transform -1 0 5980 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _48_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5428 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _49_
timestamp 1688980957
transform 1 0 4692 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _50_
timestamp 1688980957
transform 1 0 3496 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _51_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4784 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _52_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4508 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _53_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4876 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _54_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9108 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _55_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8372 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _56_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9936 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _57_
timestamp 1688980957
transform 1 0 10396 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _58_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12696 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1688980957
transform 1 0 13524 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _60_
timestamp 1688980957
transform 1 0 13984 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _61_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9844 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _62_
timestamp 1688980957
transform -1 0 8188 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _63_
timestamp 1688980957
transform -1 0 7728 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _64_
timestamp 1688980957
transform 1 0 7728 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _65_
timestamp 1688980957
transform -1 0 12420 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _66__8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11868 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _66_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11408 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11868 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1688980957
transform -1 0 7636 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1688980957
transform 1 0 10948 0 -1 13600
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1688980957
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14628 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_157
timestamp 1688980957
transform 1 0 14996 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_149 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14260 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_157
timestamp 1688980957
transform 1 0 14996 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_153
timestamp 1688980957
transform 1 0 14628 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_157
timestamp 1688980957
transform 1 0 14996 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14260 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_157
timestamp 1688980957
transform 1 0 14996 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_153
timestamp 1688980957
transform 1 0 14628 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_157
timestamp 1688980957
transform 1 0 14996 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14260 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_157
timestamp 1688980957
transform 1 0 14996 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_153
timestamp 1688980957
transform 1 0 14628 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_157
timestamp 1688980957
transform 1 0 14996 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_119
timestamp 1688980957
transform 1 0 11500 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_131
timestamp 1688980957
transform 1 0 12604 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_143
timestamp 1688980957
transform 1 0 13708 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_155
timestamp 1688980957
transform 1 0 14812 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_153
timestamp 1688980957
transform 1 0 14628 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_157
timestamp 1688980957
transform 1 0 14996 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12052 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14260 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_157
timestamp 1688980957
transform 1 0 14996 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_153
timestamp 1688980957
transform 1 0 14628 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_157
timestamp 1688980957
transform 1 0 14996 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10212 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 10948 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13156 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14260 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_157
timestamp 1688980957
transform 1 0 14996 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 9476 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 10580 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 12788 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_153
timestamp 1688980957
transform 1 0 14628 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_157
timestamp 1688980957
transform 1 0 14996 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10212 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 10948 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12052 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_149
timestamp 1688980957
transform 1 0 14260 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_157
timestamp 1688980957
transform 1 0 14996 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8372 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 10580 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 12788 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_153
timestamp 1688980957
transform 1 0 14628 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_157
timestamp 1688980957
transform 1 0 14996 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10212 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12052 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14260 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_157
timestamp 1688980957
transform 1 0 14996 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 7636 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 9476 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1688980957
transform 1 0 10580 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1688980957
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1688980957
transform 1 0 12788 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_153
timestamp 1688980957
transform 1 0 14628 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_157
timestamp 1688980957
transform 1 0 14996 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8004 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10212 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 10948 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12052 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1688980957
transform 1 0 13156 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_149
timestamp 1688980957
transform 1 0 14260 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_157
timestamp 1688980957
transform 1 0 14996 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1688980957
transform 1 0 6532 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 9476 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1688980957
transform 1 0 10580 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1688980957
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1688980957
transform 1 0 12788 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_153
timestamp 1688980957
transform 1 0 14628 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_157
timestamp 1688980957
transform 1 0 14996 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 5796 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1688980957
transform 1 0 8004 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1688980957
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1688980957
transform 1 0 10212 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1688980957
transform 1 0 10948 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12052 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1688980957
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_149
timestamp 1688980957
transform 1 0 14260 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_157
timestamp 1688980957
transform 1 0 14996 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1688980957
transform 1 0 6532 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 7636 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8372 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 9476 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1688980957
transform 1 0 10580 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1688980957
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1688980957
transform 1 0 12788 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_153
timestamp 1688980957
transform 1 0 14628 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_157
timestamp 1688980957
transform 1 0 14996 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4140 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 1688980957
transform 1 0 5428 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_57
timestamp 1688980957
transform 1 0 5796 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_65
timestamp 1688980957
transform 1 0 6532 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_73
timestamp 1688980957
transform 1 0 7268 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_85
timestamp 1688980957
transform 1 0 8372 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_97
timestamp 1688980957
transform 1 0 9476 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_109
timestamp 1688980957
transform 1 0 10580 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 10948 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12052 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13156 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_149
timestamp 1688980957
transform 1 0 14260 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_156 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14904 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4324 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_45
timestamp 1688980957
transform 1 0 4692 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_59
timestamp 1688980957
transform 1 0 5980 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_101
timestamp 1688980957
transform 1 0 9844 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_129
timestamp 1688980957
transform 1 0 12420 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_137
timestamp 1688980957
transform 1 0 13156 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1688980957
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_153
timestamp 1688980957
transform 1 0 14628 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_157
timestamp 1688980957
transform 1 0 14996 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4140 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1688980957
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_80
timestamp 1688980957
transform 1 0 7912 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_92
timestamp 1688980957
transform 1 0 9016 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_100
timestamp 1688980957
transform 1 0 9752 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 1688980957
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_133
timestamp 1688980957
transform 1 0 12788 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_145
timestamp 1688980957
transform 1 0 13892 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_157
timestamp 1688980957
transform 1 0 14996 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3220 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_37
timestamp 1688980957
transform 1 0 3956 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_46
timestamp 1688980957
transform 1 0 4784 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_54
timestamp 1688980957
transform 1 0 5520 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_63
timestamp 1688980957
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_69
timestamp 1688980957
transform 1 0 6900 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1688980957
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_100
timestamp 1688980957
transform 1 0 9752 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1688980957
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_144
timestamp 1688980957
transform 1 0 13800 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_156
timestamp 1688980957
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3036 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_31
timestamp 1688980957
transform 1 0 3404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_47
timestamp 1688980957
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_61
timestamp 1688980957
transform 1 0 6164 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_106
timestamp 1688980957
transform 1 0 10304 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_113
timestamp 1688980957
transform 1 0 10948 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_117
timestamp 1688980957
transform 1 0 11316 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_149
timestamp 1688980957
transform 1 0 14260 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_157
timestamp 1688980957
transform 1 0 14996 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_3
timestamp 1688980957
transform 1 0 828 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_7
timestamp 1688980957
transform 1 0 1196 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_11
timestamp 1688980957
transform 1 0 1564 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_23
timestamp 1688980957
transform 1 0 2668 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_33
timestamp 1688980957
transform 1 0 3588 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_43
timestamp 1688980957
transform 1 0 4508 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_49
timestamp 1688980957
transform 1 0 5060 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_57
timestamp 1688980957
transform 1 0 5796 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_75
timestamp 1688980957
transform 1 0 7452 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_97
timestamp 1688980957
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_107
timestamp 1688980957
transform 1 0 10396 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_111
timestamp 1688980957
transform 1 0 10764 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_126
timestamp 1688980957
transform 1 0 12144 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_137
timestamp 1688980957
transform 1 0 13156 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_153
timestamp 1688980957
transform 1 0 14628 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_157
timestamp 1688980957
transform 1 0 14996 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8464 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 7176 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 6992 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 9660 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 13984 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10948 0 1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform -1 0 8832 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 7452 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3220 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 1288 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 13156 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 15364 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 15364 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 15364 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 15364 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 15364 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 15364 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 15364 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 15364 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 15364 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 15364 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 15364 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 15364 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 15364 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 15364 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 15364 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 15364 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 15364 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 15364 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 15364 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 15364 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 15364 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 15364 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 15364 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 15364 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 15364 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 15364 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 15364 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 5704 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 10856 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 13432 0 1 14688
box -38 -48 130 592
<< labels >>
rlabel metal2 s 8036 14688 8036 14688 4 VGND
rlabel metal1 s 7958 15232 7958 15232 4 VPWR
rlabel metal1 s 13531 14518 13531 14518 4 _00_
rlabel metal1 s 9384 12410 9384 12410 4 _01_
rlabel metal2 s 7870 12682 7870 12682 4 _02_
rlabel metal1 s 6946 13906 6946 13906 4 _03_
rlabel metal2 s 8418 14246 8418 14246 4 _04_
rlabel metal2 s 13294 13192 13294 13192 4 _05_
rlabel metal1 s 14214 12274 14214 12274 4 _06_
rlabel metal2 s 11408 6900 11408 6900 4 _07_
rlabel metal1 s 5244 13362 5244 13362 4 _08_
rlabel metal1 s 6302 13974 6302 13974 4 _09_
rlabel metal1 s 5566 14042 5566 14042 4 _10_
rlabel metal1 s 5566 14518 5566 14518 4 _11_
rlabel metal2 s 5658 14586 5658 14586 4 _12_
rlabel metal1 s 9384 12274 9384 12274 4 _13_
rlabel metal1 s 6854 12750 6854 12750 4 _14_
rlabel metal1 s 7084 12410 7084 12410 4 _15_
rlabel metal2 s 7314 12444 7314 12444 4 _16_
rlabel metal1 s 9430 13872 9430 13872 4 _17_
rlabel metal1 s 5336 12954 5336 12954 4 _18_
rlabel metal2 s 4830 13090 4830 13090 4 _19_
rlabel metal1 s 4692 13498 4692 13498 4 _20_
rlabel metal1 s 4094 14484 4094 14484 4 _21_
rlabel metal1 s 4646 14042 4646 14042 4 _22_
rlabel metal2 s 4462 14620 4462 14620 4 _23_
rlabel metal1 s 8786 13838 8786 13838 4 _24_
rlabel metal1 s 8602 13872 8602 13872 4 _25_
rlabel metal1 s 12926 13804 12926 13804 4 _26_
rlabel metal1 s 11224 13294 11224 13294 4 _27_
rlabel metal1 s 13478 13838 13478 13838 4 _28_
rlabel metal2 s 14766 14834 14766 14834 4 clk
rlabel metal1 s 10212 13702 10212 13702 4 clknet_0_clk
rlabel metal1 s 7636 12750 7636 12750 4 clknet_1_0__leaf_clk
rlabel metal1 s 11086 12750 11086 12750 4 clknet_1_1__leaf_clk
rlabel metal1 s 5520 12070 5520 12070 4 divider\[0\]
rlabel metal2 s 6762 13328 6762 13328 4 divider\[1\]
rlabel metal1 s 5796 14382 5796 14382 4 divider\[2\]
rlabel metal2 s 10994 15351 10994 15351 4 ext_lo_en
rlabel metal1 s 8694 14926 8694 14926 4 ext_lo_n
rlabel metal1 s 7176 14926 7176 14926 4 ext_lo_p
rlabel metal1 s 9660 14586 9660 14586 4 int_lo_n
rlabel metal1 s 11454 13362 11454 13362 4 int_lo_p
rlabel metal1 s 5152 14926 5152 14926 4 int_lo_settings[0]
rlabel metal1 s 3266 14926 3266 14926 4 int_lo_settings[1]
rlabel metal1 s 1288 14926 1288 14926 4 int_lo_settings[2]
rlabel metal3 s 15234 11764 15234 11764 4 lo_n
rlabel metal3 s 13409 4148 13409 4148 4 lo_p
rlabel metal1 s 12880 14926 12880 14926 4 n_rst
rlabel metal2 s 12466 14416 12466 14416 4 net1
rlabel metal1 s 6440 14926 6440 14926 4 net10
rlabel metal1 s 7636 14042 7636 14042 4 net11
rlabel metal1 s 10304 14450 10304 14450 4 net12
rlabel metal1 s 13018 13872 13018 13872 4 net13
rlabel metal1 s 9154 14586 9154 14586 4 net2
rlabel metal1 s 12190 13906 12190 13906 4 net3
rlabel metal1 s 4830 12274 4830 12274 4 net4
rlabel metal2 s 5382 14331 5382 14331 4 net5
rlabel metal1 s 1518 14518 1518 14518 4 net6
rlabel metal1 s 13570 14450 13570 14450 4 net7
rlabel metal1 s 11776 14382 11776 14382 4 net8
rlabel metal1 s 8694 12410 8694 12410 4 net9
rlabel metal1 s 13524 14382 13524 14382 4 rst
flabel metal4 s 15200 496 15520 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 11498 496 11818 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7796 496 8116 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4094 496 4414 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 13349 496 13669 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 9647 496 9967 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 5945 496 6265 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2243 496 2563 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 14738 15600 14794 16000 0 FreeSans 280 90 0 0 clk
port 3 nsew
flabel metal2 s 10874 15600 10930 16000 0 FreeSans 280 90 0 0 ext_lo_en
port 4 nsew
flabel metal2 s 8942 15600 8998 16000 0 FreeSans 280 90 0 0 ext_lo_n
port 5 nsew
flabel metal2 s 7010 15600 7066 16000 0 FreeSans 280 90 0 0 ext_lo_p
port 6 nsew
flabel metal2 s 5078 15600 5134 16000 0 FreeSans 280 90 0 0 int_lo_settings[0]
port 7 nsew
flabel metal2 s 3146 15600 3202 16000 0 FreeSans 280 90 0 0 int_lo_settings[1]
port 8 nsew
flabel metal2 s 1214 15600 1270 16000 0 FreeSans 280 90 0 0 int_lo_settings[2]
port 9 nsew
flabel metal3 s 15600 11704 16000 11824 0 FreeSans 600 0 0 0 lo_n
port 10 nsew
flabel metal3 s 15600 3816 16000 3936 0 FreeSans 600 0 0 0 lo_p
port 11 nsew
flabel metal2 s 12806 15600 12862 16000 0 FreeSans 280 90 0 0 n_rst
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 16000 16000
string GDS_END 457902
string GDS_FILE ../gds/mixer_control.gds
string GDS_START 208040
<< end >>
