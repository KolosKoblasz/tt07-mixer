magic
tech sky130A
magscale 1 2
timestamp 1716477521
<< pwell >>
rect -1565 -761 1565 761
<< psubdiff >>
rect -1529 691 -1433 725
rect 1433 691 1529 725
rect -1529 629 -1495 691
rect 1495 629 1529 691
rect -1529 -691 -1495 -629
rect 1495 -691 1529 -629
rect -1529 -725 -1433 -691
rect 1433 -725 1529 -691
<< psubdiffcont >>
rect -1433 691 1433 725
rect -1529 -629 -1495 629
rect 1495 -629 1529 629
rect -1433 -725 1433 -691
<< poly >>
rect -1399 579 -1299 595
rect -1399 545 -1383 579
rect -1315 545 -1299 579
rect -1399 165 -1299 545
rect -1399 -545 -1299 -165
rect -1399 -579 -1383 -545
rect -1315 -579 -1299 -545
rect -1399 -595 -1299 -579
rect -1257 579 -1157 595
rect -1257 545 -1241 579
rect -1173 545 -1157 579
rect -1257 165 -1157 545
rect -1257 -545 -1157 -165
rect -1257 -579 -1241 -545
rect -1173 -579 -1157 -545
rect -1257 -595 -1157 -579
rect -1115 579 -1015 595
rect -1115 545 -1099 579
rect -1031 545 -1015 579
rect -1115 165 -1015 545
rect -1115 -545 -1015 -165
rect -1115 -579 -1099 -545
rect -1031 -579 -1015 -545
rect -1115 -595 -1015 -579
rect -973 579 -873 595
rect -973 545 -957 579
rect -889 545 -873 579
rect -973 165 -873 545
rect -973 -545 -873 -165
rect -973 -579 -957 -545
rect -889 -579 -873 -545
rect -973 -595 -873 -579
rect -831 579 -731 595
rect -831 545 -815 579
rect -747 545 -731 579
rect -831 165 -731 545
rect -831 -545 -731 -165
rect -831 -579 -815 -545
rect -747 -579 -731 -545
rect -831 -595 -731 -579
rect -689 579 -589 595
rect -689 545 -673 579
rect -605 545 -589 579
rect -689 165 -589 545
rect -689 -545 -589 -165
rect -689 -579 -673 -545
rect -605 -579 -589 -545
rect -689 -595 -589 -579
rect -547 579 -447 595
rect -547 545 -531 579
rect -463 545 -447 579
rect -547 165 -447 545
rect -547 -545 -447 -165
rect -547 -579 -531 -545
rect -463 -579 -447 -545
rect -547 -595 -447 -579
rect -405 579 -305 595
rect -405 545 -389 579
rect -321 545 -305 579
rect -405 165 -305 545
rect -405 -545 -305 -165
rect -405 -579 -389 -545
rect -321 -579 -305 -545
rect -405 -595 -305 -579
rect -263 579 -163 595
rect -263 545 -247 579
rect -179 545 -163 579
rect -263 165 -163 545
rect -263 -545 -163 -165
rect -263 -579 -247 -545
rect -179 -579 -163 -545
rect -263 -595 -163 -579
rect -121 579 -21 595
rect -121 545 -105 579
rect -37 545 -21 579
rect -121 165 -21 545
rect -121 -545 -21 -165
rect -121 -579 -105 -545
rect -37 -579 -21 -545
rect -121 -595 -21 -579
rect 21 579 121 595
rect 21 545 37 579
rect 105 545 121 579
rect 21 165 121 545
rect 21 -545 121 -165
rect 21 -579 37 -545
rect 105 -579 121 -545
rect 21 -595 121 -579
rect 163 579 263 595
rect 163 545 179 579
rect 247 545 263 579
rect 163 165 263 545
rect 163 -545 263 -165
rect 163 -579 179 -545
rect 247 -579 263 -545
rect 163 -595 263 -579
rect 305 579 405 595
rect 305 545 321 579
rect 389 545 405 579
rect 305 165 405 545
rect 305 -545 405 -165
rect 305 -579 321 -545
rect 389 -579 405 -545
rect 305 -595 405 -579
rect 447 579 547 595
rect 447 545 463 579
rect 531 545 547 579
rect 447 165 547 545
rect 447 -545 547 -165
rect 447 -579 463 -545
rect 531 -579 547 -545
rect 447 -595 547 -579
rect 589 579 689 595
rect 589 545 605 579
rect 673 545 689 579
rect 589 165 689 545
rect 589 -545 689 -165
rect 589 -579 605 -545
rect 673 -579 689 -545
rect 589 -595 689 -579
rect 731 579 831 595
rect 731 545 747 579
rect 815 545 831 579
rect 731 165 831 545
rect 731 -545 831 -165
rect 731 -579 747 -545
rect 815 -579 831 -545
rect 731 -595 831 -579
rect 873 579 973 595
rect 873 545 889 579
rect 957 545 973 579
rect 873 165 973 545
rect 873 -545 973 -165
rect 873 -579 889 -545
rect 957 -579 973 -545
rect 873 -595 973 -579
rect 1015 579 1115 595
rect 1015 545 1031 579
rect 1099 545 1115 579
rect 1015 165 1115 545
rect 1015 -545 1115 -165
rect 1015 -579 1031 -545
rect 1099 -579 1115 -545
rect 1015 -595 1115 -579
rect 1157 579 1257 595
rect 1157 545 1173 579
rect 1241 545 1257 579
rect 1157 165 1257 545
rect 1157 -545 1257 -165
rect 1157 -579 1173 -545
rect 1241 -579 1257 -545
rect 1157 -595 1257 -579
rect 1299 579 1399 595
rect 1299 545 1315 579
rect 1383 545 1399 579
rect 1299 165 1399 545
rect 1299 -545 1399 -165
rect 1299 -579 1315 -545
rect 1383 -579 1399 -545
rect 1299 -595 1399 -579
<< polycont >>
rect -1383 545 -1315 579
rect -1383 -579 -1315 -545
rect -1241 545 -1173 579
rect -1241 -579 -1173 -545
rect -1099 545 -1031 579
rect -1099 -579 -1031 -545
rect -957 545 -889 579
rect -957 -579 -889 -545
rect -815 545 -747 579
rect -815 -579 -747 -545
rect -673 545 -605 579
rect -673 -579 -605 -545
rect -531 545 -463 579
rect -531 -579 -463 -545
rect -389 545 -321 579
rect -389 -579 -321 -545
rect -247 545 -179 579
rect -247 -579 -179 -545
rect -105 545 -37 579
rect -105 -579 -37 -545
rect 37 545 105 579
rect 37 -579 105 -545
rect 179 545 247 579
rect 179 -579 247 -545
rect 321 545 389 579
rect 321 -579 389 -545
rect 463 545 531 579
rect 463 -579 531 -545
rect 605 545 673 579
rect 605 -579 673 -545
rect 747 545 815 579
rect 747 -579 815 -545
rect 889 545 957 579
rect 889 -579 957 -545
rect 1031 545 1099 579
rect 1031 -579 1099 -545
rect 1173 545 1241 579
rect 1173 -579 1241 -545
rect 1315 545 1383 579
rect 1315 -579 1383 -545
<< npolyres >>
rect -1399 -165 -1299 165
rect -1257 -165 -1157 165
rect -1115 -165 -1015 165
rect -973 -165 -873 165
rect -831 -165 -731 165
rect -689 -165 -589 165
rect -547 -165 -447 165
rect -405 -165 -305 165
rect -263 -165 -163 165
rect -121 -165 -21 165
rect 21 -165 121 165
rect 163 -165 263 165
rect 305 -165 405 165
rect 447 -165 547 165
rect 589 -165 689 165
rect 731 -165 831 165
rect 873 -165 973 165
rect 1015 -165 1115 165
rect 1157 -165 1257 165
rect 1299 -165 1399 165
<< locali >>
rect -1529 691 -1433 725
rect 1433 691 1529 725
rect -1529 629 -1495 691
rect 1495 629 1529 691
rect -1399 545 -1383 579
rect -1315 545 -1299 579
rect -1257 545 -1241 579
rect -1173 545 -1157 579
rect -1115 545 -1099 579
rect -1031 545 -1015 579
rect -973 545 -957 579
rect -889 545 -873 579
rect -831 545 -815 579
rect -747 545 -731 579
rect -689 545 -673 579
rect -605 545 -589 579
rect -547 545 -531 579
rect -463 545 -447 579
rect -405 545 -389 579
rect -321 545 -305 579
rect -263 545 -247 579
rect -179 545 -163 579
rect -121 545 -105 579
rect -37 545 -21 579
rect 21 545 37 579
rect 105 545 121 579
rect 163 545 179 579
rect 247 545 263 579
rect 305 545 321 579
rect 389 545 405 579
rect 447 545 463 579
rect 531 545 547 579
rect 589 545 605 579
rect 673 545 689 579
rect 731 545 747 579
rect 815 545 831 579
rect 873 545 889 579
rect 957 545 973 579
rect 1015 545 1031 579
rect 1099 545 1115 579
rect 1157 545 1173 579
rect 1241 545 1257 579
rect 1299 545 1315 579
rect 1383 545 1399 579
rect -1399 -579 -1383 -545
rect -1315 -579 -1299 -545
rect -1257 -579 -1241 -545
rect -1173 -579 -1157 -545
rect -1115 -579 -1099 -545
rect -1031 -579 -1015 -545
rect -973 -579 -957 -545
rect -889 -579 -873 -545
rect -831 -579 -815 -545
rect -747 -579 -731 -545
rect -689 -579 -673 -545
rect -605 -579 -589 -545
rect -547 -579 -531 -545
rect -463 -579 -447 -545
rect -405 -579 -389 -545
rect -321 -579 -305 -545
rect -263 -579 -247 -545
rect -179 -579 -163 -545
rect -121 -579 -105 -545
rect -37 -579 -21 -545
rect 21 -579 37 -545
rect 105 -579 121 -545
rect 163 -579 179 -545
rect 247 -579 263 -545
rect 305 -579 321 -545
rect 389 -579 405 -545
rect 447 -579 463 -545
rect 531 -579 547 -545
rect 589 -579 605 -545
rect 673 -579 689 -545
rect 731 -579 747 -545
rect 815 -579 831 -545
rect 873 -579 889 -545
rect 957 -579 973 -545
rect 1015 -579 1031 -545
rect 1099 -579 1115 -545
rect 1157 -579 1173 -545
rect 1241 -579 1257 -545
rect 1299 -579 1315 -545
rect 1383 -579 1399 -545
rect -1529 -691 -1495 -629
rect 1495 -691 1529 -629
rect -1529 -725 -1433 -691
rect 1433 -725 1529 -691
<< viali >>
rect -1383 545 -1315 579
rect -1241 545 -1173 579
rect -1099 545 -1031 579
rect -957 545 -889 579
rect -815 545 -747 579
rect -673 545 -605 579
rect -531 545 -463 579
rect -389 545 -321 579
rect -247 545 -179 579
rect -105 545 -37 579
rect 37 545 105 579
rect 179 545 247 579
rect 321 545 389 579
rect 463 545 531 579
rect 605 545 673 579
rect 747 545 815 579
rect 889 545 957 579
rect 1031 545 1099 579
rect 1173 545 1241 579
rect 1315 545 1383 579
rect -1383 182 -1315 545
rect -1241 182 -1173 545
rect -1099 182 -1031 545
rect -957 182 -889 545
rect -815 182 -747 545
rect -673 182 -605 545
rect -531 182 -463 545
rect -389 182 -321 545
rect -247 182 -179 545
rect -105 182 -37 545
rect 37 182 105 545
rect 179 182 247 545
rect 321 182 389 545
rect 463 182 531 545
rect 605 182 673 545
rect 747 182 815 545
rect 889 182 957 545
rect 1031 182 1099 545
rect 1173 182 1241 545
rect 1315 182 1383 545
rect -1383 -545 -1315 -182
rect -1241 -545 -1173 -182
rect -1099 -545 -1031 -182
rect -957 -545 -889 -182
rect -815 -545 -747 -182
rect -673 -545 -605 -182
rect -531 -545 -463 -182
rect -389 -545 -321 -182
rect -247 -545 -179 -182
rect -105 -545 -37 -182
rect 37 -545 105 -182
rect 179 -545 247 -182
rect 321 -545 389 -182
rect 463 -545 531 -182
rect 605 -545 673 -182
rect 747 -545 815 -182
rect 889 -545 957 -182
rect 1031 -545 1099 -182
rect 1173 -545 1241 -182
rect 1315 -545 1383 -182
rect -1383 -579 -1315 -545
rect -1241 -579 -1173 -545
rect -1099 -579 -1031 -545
rect -957 -579 -889 -545
rect -815 -579 -747 -545
rect -673 -579 -605 -545
rect -531 -579 -463 -545
rect -389 -579 -321 -545
rect -247 -579 -179 -545
rect -105 -579 -37 -545
rect 37 -579 105 -545
rect 179 -579 247 -545
rect 321 -579 389 -545
rect 463 -579 531 -545
rect 605 -579 673 -545
rect 747 -579 815 -545
rect 889 -579 957 -545
rect 1031 -579 1099 -545
rect 1173 -579 1241 -545
rect 1315 -579 1383 -545
<< metal1 >>
rect -1389 579 -1309 591
rect -1389 182 -1383 579
rect -1315 182 -1309 579
rect -1389 170 -1309 182
rect -1247 579 -1167 591
rect -1247 182 -1241 579
rect -1173 182 -1167 579
rect -1247 170 -1167 182
rect -1105 579 -1025 591
rect -1105 182 -1099 579
rect -1031 182 -1025 579
rect -1105 170 -1025 182
rect -963 579 -883 591
rect -963 182 -957 579
rect -889 182 -883 579
rect -963 170 -883 182
rect -821 579 -741 591
rect -821 182 -815 579
rect -747 182 -741 579
rect -821 170 -741 182
rect -679 579 -599 591
rect -679 182 -673 579
rect -605 182 -599 579
rect -679 170 -599 182
rect -537 579 -457 591
rect -537 182 -531 579
rect -463 182 -457 579
rect -537 170 -457 182
rect -395 579 -315 591
rect -395 182 -389 579
rect -321 182 -315 579
rect -395 170 -315 182
rect -253 579 -173 591
rect -253 182 -247 579
rect -179 182 -173 579
rect -253 170 -173 182
rect -111 579 -31 591
rect -111 182 -105 579
rect -37 182 -31 579
rect -111 170 -31 182
rect 31 579 111 591
rect 31 182 37 579
rect 105 182 111 579
rect 31 170 111 182
rect 173 579 253 591
rect 173 182 179 579
rect 247 182 253 579
rect 173 170 253 182
rect 315 579 395 591
rect 315 182 321 579
rect 389 182 395 579
rect 315 170 395 182
rect 457 579 537 591
rect 457 182 463 579
rect 531 182 537 579
rect 457 170 537 182
rect 599 579 679 591
rect 599 182 605 579
rect 673 182 679 579
rect 599 170 679 182
rect 741 579 821 591
rect 741 182 747 579
rect 815 182 821 579
rect 741 170 821 182
rect 883 579 963 591
rect 883 182 889 579
rect 957 182 963 579
rect 883 170 963 182
rect 1025 579 1105 591
rect 1025 182 1031 579
rect 1099 182 1105 579
rect 1025 170 1105 182
rect 1167 579 1247 591
rect 1167 182 1173 579
rect 1241 182 1247 579
rect 1167 170 1247 182
rect 1309 579 1389 591
rect 1309 182 1315 579
rect 1383 182 1389 579
rect 1309 170 1389 182
rect -1389 -182 -1309 -170
rect -1389 -579 -1383 -182
rect -1315 -579 -1309 -182
rect -1389 -591 -1309 -579
rect -1247 -182 -1167 -170
rect -1247 -579 -1241 -182
rect -1173 -579 -1167 -182
rect -1247 -591 -1167 -579
rect -1105 -182 -1025 -170
rect -1105 -579 -1099 -182
rect -1031 -579 -1025 -182
rect -1105 -591 -1025 -579
rect -963 -182 -883 -170
rect -963 -579 -957 -182
rect -889 -579 -883 -182
rect -963 -591 -883 -579
rect -821 -182 -741 -170
rect -821 -579 -815 -182
rect -747 -579 -741 -182
rect -821 -591 -741 -579
rect -679 -182 -599 -170
rect -679 -579 -673 -182
rect -605 -579 -599 -182
rect -679 -591 -599 -579
rect -537 -182 -457 -170
rect -537 -579 -531 -182
rect -463 -579 -457 -182
rect -537 -591 -457 -579
rect -395 -182 -315 -170
rect -395 -579 -389 -182
rect -321 -579 -315 -182
rect -395 -591 -315 -579
rect -253 -182 -173 -170
rect -253 -579 -247 -182
rect -179 -579 -173 -182
rect -253 -591 -173 -579
rect -111 -182 -31 -170
rect -111 -579 -105 -182
rect -37 -579 -31 -182
rect -111 -591 -31 -579
rect 31 -182 111 -170
rect 31 -579 37 -182
rect 105 -579 111 -182
rect 31 -591 111 -579
rect 173 -182 253 -170
rect 173 -579 179 -182
rect 247 -579 253 -182
rect 173 -591 253 -579
rect 315 -182 395 -170
rect 315 -579 321 -182
rect 389 -579 395 -182
rect 315 -591 395 -579
rect 457 -182 537 -170
rect 457 -579 463 -182
rect 531 -579 537 -182
rect 457 -591 537 -579
rect 599 -182 679 -170
rect 599 -579 605 -182
rect 673 -579 679 -182
rect 599 -591 679 -579
rect 741 -182 821 -170
rect 741 -579 747 -182
rect 815 -579 821 -182
rect 741 -591 821 -579
rect 883 -182 963 -170
rect 883 -579 889 -182
rect 957 -579 963 -182
rect 883 -591 963 -579
rect 1025 -182 1105 -170
rect 1025 -579 1031 -182
rect 1099 -579 1105 -182
rect 1025 -591 1105 -579
rect 1167 -182 1247 -170
rect 1167 -579 1173 -182
rect 1241 -579 1247 -182
rect 1167 -591 1247 -579
rect 1309 -182 1389 -170
rect 1309 -579 1315 -182
rect 1383 -579 1389 -182
rect 1309 -591 1389 -579
<< properties >>
string FIXED_BBOX -1512 -708 1512 708
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.5 l 1.650 m 1 nx 20 wmin 0.330 lmin 1.650 rho 48.2 val 159.06 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
