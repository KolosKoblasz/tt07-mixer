magic
tech sky130A
magscale 1 2
timestamp 1716477521
<< pwell >>
rect -361 -2702 361 2702
<< psubdiff >>
rect -325 2632 -229 2666
rect 229 2632 325 2666
rect -325 2570 -291 2632
rect 291 2570 325 2632
rect -325 -2632 -291 -2570
rect 291 -2632 325 -2570
rect -325 -2666 -229 -2632
rect 229 -2666 325 -2632
<< psubdiffcont >>
rect -229 2632 229 2666
rect -325 -2570 -291 2570
rect 291 -2570 325 2570
rect -229 -2666 229 -2632
<< poly >>
rect -195 2520 -129 2536
rect -195 2486 -179 2520
rect -145 2486 -129 2520
rect -195 2106 -129 2486
rect -195 1396 -129 1776
rect -195 1362 -179 1396
rect -145 1362 -129 1396
rect -195 1346 -129 1362
rect -87 2520 -21 2536
rect -87 2486 -71 2520
rect -37 2486 -21 2520
rect -87 2106 -21 2486
rect -87 1396 -21 1776
rect -87 1362 -71 1396
rect -37 1362 -21 1396
rect -87 1346 -21 1362
rect 21 2520 87 2536
rect 21 2486 37 2520
rect 71 2486 87 2520
rect 21 2106 87 2486
rect 21 1396 87 1776
rect 21 1362 37 1396
rect 71 1362 87 1396
rect 21 1346 87 1362
rect 129 2520 195 2536
rect 129 2486 145 2520
rect 179 2486 195 2520
rect 129 2106 195 2486
rect 129 1396 195 1776
rect 129 1362 145 1396
rect 179 1362 195 1396
rect 129 1346 195 1362
rect -195 1226 -129 1242
rect -195 1192 -179 1226
rect -145 1192 -129 1226
rect -195 812 -129 1192
rect -195 102 -129 482
rect -195 68 -179 102
rect -145 68 -129 102
rect -195 52 -129 68
rect -87 1226 -21 1242
rect -87 1192 -71 1226
rect -37 1192 -21 1226
rect -87 812 -21 1192
rect -87 102 -21 482
rect -87 68 -71 102
rect -37 68 -21 102
rect -87 52 -21 68
rect 21 1226 87 1242
rect 21 1192 37 1226
rect 71 1192 87 1226
rect 21 812 87 1192
rect 21 102 87 482
rect 21 68 37 102
rect 71 68 87 102
rect 21 52 87 68
rect 129 1226 195 1242
rect 129 1192 145 1226
rect 179 1192 195 1226
rect 129 812 195 1192
rect 129 102 195 482
rect 129 68 145 102
rect 179 68 195 102
rect 129 52 195 68
rect -195 -68 -129 -52
rect -195 -102 -179 -68
rect -145 -102 -129 -68
rect -195 -482 -129 -102
rect -195 -1192 -129 -812
rect -195 -1226 -179 -1192
rect -145 -1226 -129 -1192
rect -195 -1242 -129 -1226
rect -87 -68 -21 -52
rect -87 -102 -71 -68
rect -37 -102 -21 -68
rect -87 -482 -21 -102
rect -87 -1192 -21 -812
rect -87 -1226 -71 -1192
rect -37 -1226 -21 -1192
rect -87 -1242 -21 -1226
rect 21 -68 87 -52
rect 21 -102 37 -68
rect 71 -102 87 -68
rect 21 -482 87 -102
rect 21 -1192 87 -812
rect 21 -1226 37 -1192
rect 71 -1226 87 -1192
rect 21 -1242 87 -1226
rect 129 -68 195 -52
rect 129 -102 145 -68
rect 179 -102 195 -68
rect 129 -482 195 -102
rect 129 -1192 195 -812
rect 129 -1226 145 -1192
rect 179 -1226 195 -1192
rect 129 -1242 195 -1226
rect -195 -1362 -129 -1346
rect -195 -1396 -179 -1362
rect -145 -1396 -129 -1362
rect -195 -1776 -129 -1396
rect -195 -2486 -129 -2106
rect -195 -2520 -179 -2486
rect -145 -2520 -129 -2486
rect -195 -2536 -129 -2520
rect -87 -1362 -21 -1346
rect -87 -1396 -71 -1362
rect -37 -1396 -21 -1362
rect -87 -1776 -21 -1396
rect -87 -2486 -21 -2106
rect -87 -2520 -71 -2486
rect -37 -2520 -21 -2486
rect -87 -2536 -21 -2520
rect 21 -1362 87 -1346
rect 21 -1396 37 -1362
rect 71 -1396 87 -1362
rect 21 -1776 87 -1396
rect 21 -2486 87 -2106
rect 21 -2520 37 -2486
rect 71 -2520 87 -2486
rect 21 -2536 87 -2520
rect 129 -1362 195 -1346
rect 129 -1396 145 -1362
rect 179 -1396 195 -1362
rect 129 -1776 195 -1396
rect 129 -2486 195 -2106
rect 129 -2520 145 -2486
rect 179 -2520 195 -2486
rect 129 -2536 195 -2520
<< polycont >>
rect -179 2486 -145 2520
rect -179 1362 -145 1396
rect -71 2486 -37 2520
rect -71 1362 -37 1396
rect 37 2486 71 2520
rect 37 1362 71 1396
rect 145 2486 179 2520
rect 145 1362 179 1396
rect -179 1192 -145 1226
rect -179 68 -145 102
rect -71 1192 -37 1226
rect -71 68 -37 102
rect 37 1192 71 1226
rect 37 68 71 102
rect 145 1192 179 1226
rect 145 68 179 102
rect -179 -102 -145 -68
rect -179 -1226 -145 -1192
rect -71 -102 -37 -68
rect -71 -1226 -37 -1192
rect 37 -102 71 -68
rect 37 -1226 71 -1192
rect 145 -102 179 -68
rect 145 -1226 179 -1192
rect -179 -1396 -145 -1362
rect -179 -2520 -145 -2486
rect -71 -1396 -37 -1362
rect -71 -2520 -37 -2486
rect 37 -1396 71 -1362
rect 37 -2520 71 -2486
rect 145 -1396 179 -1362
rect 145 -2520 179 -2486
<< npolyres >>
rect -195 1776 -129 2106
rect -87 1776 -21 2106
rect 21 1776 87 2106
rect 129 1776 195 2106
rect -195 482 -129 812
rect -87 482 -21 812
rect 21 482 87 812
rect 129 482 195 812
rect -195 -812 -129 -482
rect -87 -812 -21 -482
rect 21 -812 87 -482
rect 129 -812 195 -482
rect -195 -2106 -129 -1776
rect -87 -2106 -21 -1776
rect 21 -2106 87 -1776
rect 129 -2106 195 -1776
<< locali >>
rect -325 2632 -229 2666
rect 229 2632 325 2666
rect -325 2570 -291 2632
rect 291 2570 325 2632
rect -195 2486 -179 2520
rect -145 2486 -129 2520
rect -87 2486 -71 2520
rect -37 2486 -21 2520
rect 21 2486 37 2520
rect 71 2486 87 2520
rect 129 2486 145 2520
rect 179 2486 195 2520
rect -195 1362 -179 1396
rect -145 1362 -129 1396
rect -87 1362 -71 1396
rect -37 1362 -21 1396
rect 21 1362 37 1396
rect 71 1362 87 1396
rect 129 1362 145 1396
rect 179 1362 195 1396
rect -195 1192 -179 1226
rect -145 1192 -129 1226
rect -87 1192 -71 1226
rect -37 1192 -21 1226
rect 21 1192 37 1226
rect 71 1192 87 1226
rect 129 1192 145 1226
rect 179 1192 195 1226
rect -195 68 -179 102
rect -145 68 -129 102
rect -87 68 -71 102
rect -37 68 -21 102
rect 21 68 37 102
rect 71 68 87 102
rect 129 68 145 102
rect 179 68 195 102
rect -195 -102 -179 -68
rect -145 -102 -129 -68
rect -87 -102 -71 -68
rect -37 -102 -21 -68
rect 21 -102 37 -68
rect 71 -102 87 -68
rect 129 -102 145 -68
rect 179 -102 195 -68
rect -195 -1226 -179 -1192
rect -145 -1226 -129 -1192
rect -87 -1226 -71 -1192
rect -37 -1226 -21 -1192
rect 21 -1226 37 -1192
rect 71 -1226 87 -1192
rect 129 -1226 145 -1192
rect 179 -1226 195 -1192
rect -195 -1396 -179 -1362
rect -145 -1396 -129 -1362
rect -87 -1396 -71 -1362
rect -37 -1396 -21 -1362
rect 21 -1396 37 -1362
rect 71 -1396 87 -1362
rect 129 -1396 145 -1362
rect 179 -1396 195 -1362
rect -195 -2520 -179 -2486
rect -145 -2520 -129 -2486
rect -87 -2520 -71 -2486
rect -37 -2520 -21 -2486
rect 21 -2520 37 -2486
rect 71 -2520 87 -2486
rect 129 -2520 145 -2486
rect 179 -2520 195 -2486
rect -325 -2632 -291 -2570
rect 291 -2632 325 -2570
rect -325 -2666 -229 -2632
rect 229 -2666 325 -2632
<< viali >>
rect -179 2486 -145 2520
rect -71 2486 -37 2520
rect 37 2486 71 2520
rect 145 2486 179 2520
rect -179 2123 -145 2486
rect -71 2123 -37 2486
rect 37 2123 71 2486
rect 145 2123 179 2486
rect -179 1396 -145 1759
rect -71 1396 -37 1759
rect 37 1396 71 1759
rect 145 1396 179 1759
rect -179 1362 -145 1396
rect -71 1362 -37 1396
rect 37 1362 71 1396
rect 145 1362 179 1396
rect -179 1192 -145 1226
rect -71 1192 -37 1226
rect 37 1192 71 1226
rect 145 1192 179 1226
rect -179 829 -145 1192
rect -71 829 -37 1192
rect 37 829 71 1192
rect 145 829 179 1192
rect -179 102 -145 465
rect -71 102 -37 465
rect 37 102 71 465
rect 145 102 179 465
rect -179 68 -145 102
rect -71 68 -37 102
rect 37 68 71 102
rect 145 68 179 102
rect -179 -102 -145 -68
rect -71 -102 -37 -68
rect 37 -102 71 -68
rect 145 -102 179 -68
rect -179 -465 -145 -102
rect -71 -465 -37 -102
rect 37 -465 71 -102
rect 145 -465 179 -102
rect -179 -1192 -145 -829
rect -71 -1192 -37 -829
rect 37 -1192 71 -829
rect 145 -1192 179 -829
rect -179 -1226 -145 -1192
rect -71 -1226 -37 -1192
rect 37 -1226 71 -1192
rect 145 -1226 179 -1192
rect -179 -1396 -145 -1362
rect -71 -1396 -37 -1362
rect 37 -1396 71 -1362
rect 145 -1396 179 -1362
rect -179 -1759 -145 -1396
rect -71 -1759 -37 -1396
rect 37 -1759 71 -1396
rect 145 -1759 179 -1396
rect -179 -2486 -145 -2123
rect -71 -2486 -37 -2123
rect 37 -2486 71 -2123
rect 145 -2486 179 -2123
rect -179 -2520 -145 -2486
rect -71 -2520 -37 -2486
rect 37 -2520 71 -2486
rect 145 -2520 179 -2486
<< metal1 >>
rect -185 2520 -139 2532
rect -185 2123 -179 2520
rect -145 2123 -139 2520
rect -185 2111 -139 2123
rect -77 2520 -31 2532
rect -77 2123 -71 2520
rect -37 2123 -31 2520
rect -77 2111 -31 2123
rect 31 2520 77 2532
rect 31 2123 37 2520
rect 71 2123 77 2520
rect 31 2111 77 2123
rect 139 2520 185 2532
rect 139 2123 145 2520
rect 179 2123 185 2520
rect 139 2111 185 2123
rect -185 1759 -139 1771
rect -185 1362 -179 1759
rect -145 1362 -139 1759
rect -185 1350 -139 1362
rect -77 1759 -31 1771
rect -77 1362 -71 1759
rect -37 1362 -31 1759
rect -77 1350 -31 1362
rect 31 1759 77 1771
rect 31 1362 37 1759
rect 71 1362 77 1759
rect 31 1350 77 1362
rect 139 1759 185 1771
rect 139 1362 145 1759
rect 179 1362 185 1759
rect 139 1350 185 1362
rect -185 1226 -139 1238
rect -185 829 -179 1226
rect -145 829 -139 1226
rect -185 817 -139 829
rect -77 1226 -31 1238
rect -77 829 -71 1226
rect -37 829 -31 1226
rect -77 817 -31 829
rect 31 1226 77 1238
rect 31 829 37 1226
rect 71 829 77 1226
rect 31 817 77 829
rect 139 1226 185 1238
rect 139 829 145 1226
rect 179 829 185 1226
rect 139 817 185 829
rect -185 465 -139 477
rect -185 68 -179 465
rect -145 68 -139 465
rect -185 56 -139 68
rect -77 465 -31 477
rect -77 68 -71 465
rect -37 68 -31 465
rect -77 56 -31 68
rect 31 465 77 477
rect 31 68 37 465
rect 71 68 77 465
rect 31 56 77 68
rect 139 465 185 477
rect 139 68 145 465
rect 179 68 185 465
rect 139 56 185 68
rect -185 -68 -139 -56
rect -185 -465 -179 -68
rect -145 -465 -139 -68
rect -185 -477 -139 -465
rect -77 -68 -31 -56
rect -77 -465 -71 -68
rect -37 -465 -31 -68
rect -77 -477 -31 -465
rect 31 -68 77 -56
rect 31 -465 37 -68
rect 71 -465 77 -68
rect 31 -477 77 -465
rect 139 -68 185 -56
rect 139 -465 145 -68
rect 179 -465 185 -68
rect 139 -477 185 -465
rect -185 -829 -139 -817
rect -185 -1226 -179 -829
rect -145 -1226 -139 -829
rect -185 -1238 -139 -1226
rect -77 -829 -31 -817
rect -77 -1226 -71 -829
rect -37 -1226 -31 -829
rect -77 -1238 -31 -1226
rect 31 -829 77 -817
rect 31 -1226 37 -829
rect 71 -1226 77 -829
rect 31 -1238 77 -1226
rect 139 -829 185 -817
rect 139 -1226 145 -829
rect 179 -1226 185 -829
rect 139 -1238 185 -1226
rect -185 -1362 -139 -1350
rect -185 -1759 -179 -1362
rect -145 -1759 -139 -1362
rect -185 -1771 -139 -1759
rect -77 -1362 -31 -1350
rect -77 -1759 -71 -1362
rect -37 -1759 -31 -1362
rect -77 -1771 -31 -1759
rect 31 -1362 77 -1350
rect 31 -1759 37 -1362
rect 71 -1759 77 -1362
rect 31 -1771 77 -1759
rect 139 -1362 185 -1350
rect 139 -1759 145 -1362
rect 179 -1759 185 -1362
rect 139 -1771 185 -1759
rect -185 -2123 -139 -2111
rect -185 -2520 -179 -2123
rect -145 -2520 -139 -2123
rect -185 -2532 -139 -2520
rect -77 -2123 -31 -2111
rect -77 -2520 -71 -2123
rect -37 -2520 -31 -2123
rect -77 -2532 -31 -2520
rect 31 -2123 77 -2111
rect 31 -2520 37 -2123
rect 71 -2520 77 -2123
rect 31 -2532 77 -2520
rect 139 -2123 185 -2111
rect 139 -2520 145 -2123
rect 179 -2520 185 -2123
rect 139 -2532 185 -2520
<< properties >>
string FIXED_BBOX -308 -2649 308 2649
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.330 l 1.650 m 4 nx 4 wmin 0.330 lmin 1.650 rho 48.2 val 241.0 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
