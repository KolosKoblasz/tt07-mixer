magic
tech sky130A
magscale 1 2
timestamp 1716455288
<< error_p >>
rect -101 252 -33 258
rect 33 252 101 258
rect -101 218 -89 252
rect 33 218 45 252
rect -101 212 -33 218
rect 33 212 101 218
rect -101 -218 -33 -212
rect 33 -218 101 -212
rect -101 -252 -89 -218
rect 33 -252 45 -218
rect -101 -258 -33 -252
rect 33 -258 101 -252
<< pwell >>
rect -301 -390 301 390
<< nmos >>
rect -105 -180 -29 180
rect 29 -180 105 180
<< ndiff >>
rect -163 168 -105 180
rect -163 -168 -151 168
rect -117 -168 -105 168
rect -163 -180 -105 -168
rect -29 168 29 180
rect -29 -168 -17 168
rect 17 -168 29 168
rect -29 -180 29 -168
rect 105 168 163 180
rect 105 -168 117 168
rect 151 -168 163 168
rect 105 -180 163 -168
<< ndiffc >>
rect -151 -168 -117 168
rect -17 -168 17 168
rect 117 -168 151 168
<< psubdiff >>
rect -265 320 -169 354
rect 169 320 265 354
rect -265 258 -231 320
rect 231 258 265 320
rect -265 -320 -231 -258
rect 231 -320 265 -258
rect -265 -354 -169 -320
rect 169 -354 265 -320
<< psubdiffcont >>
rect -169 320 169 354
rect -265 -258 -231 258
rect 231 -258 265 258
rect -169 -354 169 -320
<< poly >>
rect -105 252 -29 268
rect -105 218 -89 252
rect -45 218 -29 252
rect -105 180 -29 218
rect 29 252 105 268
rect 29 218 45 252
rect 89 218 105 252
rect 29 180 105 218
rect -105 -218 -29 -180
rect -105 -252 -89 -218
rect -45 -252 -29 -218
rect -105 -268 -29 -252
rect 29 -218 105 -180
rect 29 -252 45 -218
rect 89 -252 105 -218
rect 29 -268 105 -252
<< polycont >>
rect -89 218 -45 252
rect 45 218 89 252
rect -89 -252 -45 -218
rect 45 -252 89 -218
<< locali >>
rect -265 320 -169 354
rect 169 320 265 354
rect -265 258 -231 320
rect 231 258 265 320
rect -105 218 -89 252
rect -45 218 -29 252
rect 29 218 45 252
rect 89 218 105 252
rect -151 168 -117 184
rect -151 -184 -117 -168
rect -17 168 17 184
rect -17 -184 17 -168
rect 117 168 151 184
rect 117 -184 151 -168
rect -105 -252 -89 -218
rect -45 -252 -29 -218
rect 29 -252 45 -218
rect 89 -252 105 -218
rect -265 -320 -231 -258
rect 231 -320 265 -258
rect -265 -354 -169 -320
rect 169 -354 265 -320
<< viali >>
rect -89 218 -45 252
rect 45 218 89 252
rect -151 -168 -117 168
rect -17 -168 17 168
rect 117 -168 151 168
rect -89 -252 -45 -218
rect 45 -252 89 -218
<< metal1 >>
rect -101 252 -33 258
rect -101 218 -89 252
rect -45 218 -33 252
rect -101 212 -33 218
rect 33 252 101 258
rect 33 218 45 252
rect 89 218 101 252
rect 33 212 101 218
rect -157 168 -111 180
rect -157 -168 -151 168
rect -117 -168 -111 168
rect -157 -180 -111 -168
rect -23 168 23 180
rect -23 -168 -17 168
rect 17 -168 23 168
rect -23 -180 23 -168
rect 111 168 157 180
rect 111 -168 117 168
rect 151 -168 157 168
rect 111 -180 157 -168
rect -101 -218 -33 -212
rect -101 -252 -89 -218
rect -45 -252 -33 -218
rect -101 -258 -33 -252
rect 33 -218 101 -212
rect 33 -252 45 -218
rect 89 -252 101 -218
rect 33 -258 101 -252
<< properties >>
string FIXED_BBOX -248 -337 248 337
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.8 l 0.38 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
